
//
// Verific Verilog Description of module test_periph_assembly
//

module test_periph_assembly (pins, sys_w_addr, sys_r_addr, sys_w_line, 
            sys_r_line, sys_w, sys_r, rst, clk);   // test_periph_assembly.v(6)
    inout [127:0]pins;   // test_periph_assembly.v(7)
    input [31:0]sys_w_addr;   // test_periph_assembly.v(10)
    input [31:0]sys_r_addr;   // test_periph_assembly.v(11)
    input [31:0]sys_w_line;   // test_periph_assembly.v(12)
    output [31:0]sys_r_line;   // test_periph_assembly.v(13)
    input sys_w;   // test_periph_assembly.v(14)
    input sys_r;   // test_periph_assembly.v(15)
    input rst;   // test_periph_assembly.v(19)
    input clk;   // test_periph_assembly.v(18)
    
    wire [31:0]g0_in;   // test_periph_assembly.v(39)
    wire [31:0]g1_in;   // test_periph_assembly.v(39)
    wire [31:0]g2_in;   // test_periph_assembly.v(39)
    wire [31:0]g3_in;   // test_periph_assembly.v(39)
    wire [31:0]mx0_f0_out;   // test_periph_assembly.v(48)
    wire [31:0]mx0_f1_out;   // test_periph_assembly.v(48)
    wire [31:0]mx0_f2_out;   // test_periph_assembly.v(48)
    wire [31:0]mx0_f3_out;   // test_periph_assembly.v(48)
    wire [31:0]mx1_f0_out;   // test_periph_assembly.v(49)
    wire [31:0]mx1_f1_out;   // test_periph_assembly.v(49)
    wire [31:0]mx1_f2_out;   // test_periph_assembly.v(49)
    wire [31:0]mx1_f3_out;   // test_periph_assembly.v(49)
    wire [31:0]mx2_f0_out;   // test_periph_assembly.v(50)
    wire [31:0]mx2_f1_out;   // test_periph_assembly.v(50)
    wire [31:0]mx2_f2_out;   // test_periph_assembly.v(50)
    wire [31:0]mx2_f3_out;   // test_periph_assembly.v(50)
    wire [31:0]mx3_f0_out;   // test_periph_assembly.v(51)
    wire [31:0]mx3_f1_out;   // test_periph_assembly.v(51)
    wire [31:0]mx3_f2_out;   // test_periph_assembly.v(51)
    wire [31:0]mx3_f3_out;   // test_periph_assembly.v(51)
    wire [31:0]mx0_f0_dir;   // test_periph_assembly.v(58)
    wire [31:0]mx0_f1_dir;   // test_periph_assembly.v(58)
    wire [31:0]mx0_f2_dir;   // test_periph_assembly.v(58)
    wire [31:0]mx0_f3_dir;   // test_periph_assembly.v(58)
    wire [31:0]mx1_f0_dir;   // test_periph_assembly.v(59)
    wire [31:0]mx1_f1_dir;   // test_periph_assembly.v(59)
    wire [31:0]mx1_f2_dir;   // test_periph_assembly.v(59)
    wire [31:0]mx1_f3_dir;   // test_periph_assembly.v(59)
    wire [31:0]mx2_f0_dir;   // test_periph_assembly.v(60)
    wire [31:0]mx2_f1_dir;   // test_periph_assembly.v(60)
    wire [31:0]mx2_f2_dir;   // test_periph_assembly.v(60)
    wire [31:0]mx2_f3_dir;   // test_periph_assembly.v(60)
    wire [31:0]mx3_f0_dir;   // test_periph_assembly.v(61)
    wire [31:0]mx3_f1_dir;   // test_periph_assembly.v(61)
    wire [31:0]mx3_f2_dir;   // test_periph_assembly.v(61)
    wire [31:0]mx3_f3_dir;   // test_periph_assembly.v(61)
    
    gpio chip0 (.gpio_out({mx0_f0_out}), .gpio_in({g0_in}), .gpio_dir({mx0_f0_dir}), 
         .addr({32'b00000000000000000000000000001010}), .sys_w_addr({sys_w_addr}), 
         .sys_r_addr({sys_r_addr}), .sys_w_line({sys_w_line}), .sys_r_line({sys_r_line}), 
         .sys_w(sys_w), .sys_r(sys_r), .rst(rst), .clk(clk));   // test_periph_assembly.v(41)
    gpio chip1 (.gpio_out({mx1_f0_out}), .gpio_in({g1_in}), .gpio_dir({mx1_f0_dir}), 
         .addr({32'b00000000000000000000000000001100}), .sys_w_addr({sys_w_addr}), 
         .sys_r_addr({sys_r_addr}), .sys_w_line({sys_w_line}), .sys_r_line({sys_r_line}), 
         .sys_w(sys_w), .sys_r(sys_r), .rst(rst), .clk(clk));   // test_periph_assembly.v(42)
    gpio chip2 (.gpio_out({mx2_f0_out}), .gpio_in({g2_in}), .gpio_dir({mx2_f0_dir}), 
         .addr({32'b00000000000000000000000000001110}), .sys_w_addr({sys_w_addr}), 
         .sys_r_addr({sys_r_addr}), .sys_w_line({sys_w_line}), .sys_r_line({sys_r_line}), 
         .sys_w(sys_w), .sys_r(sys_r), .rst(rst), .clk(clk));   // test_periph_assembly.v(43)
    gpio chip3 (.gpio_out({mx3_f0_out}), .gpio_in({g3_in}), .gpio_dir({mx3_f0_dir}), 
         .addr({32'b00000000000000000000000000010000}), .sys_w_addr({sys_w_addr}), 
         .sys_r_addr({sys_r_addr}), .sys_w_line({sys_w_line}), .sys_r_line({sys_r_line}), 
         .sys_w(sys_w), .sys_r(sys_r), .rst(rst), .clk(clk));   // test_periph_assembly.v(44)
    gpio_mux mx0 (.pins({pins[31:0]}), .func0_in({g0_in}), .func0_out({mx0_f0_out}), 
            .func1_out({mx0_f1_out}), .func2_out({mx0_f2_out}), .func3_out({mx0_f3_out}), 
            .func0_dir({mx0_f0_dir}), .func1_dir({mx0_f1_dir}), .func2_dir({mx0_f2_dir}), 
            .func3_dir({mx0_f3_dir}), .addr({32'b00000000000000000000000000000010}), 
            .sys_w_addr({sys_w_addr}), .sys_r_addr({sys_r_addr}), .sys_w_line({sys_w_line}), 
            .sys_r_line({sys_r_line}), .sys_w(sys_w), .sys_r(sys_r), .rst(rst), 
            .clk(clk));   // test_periph_assembly.v(63)
    gpio_mux mx1 (.pins({pins[63:32]}), .func0_in({g1_in}), .func0_out({mx1_f0_out}), 
            .func1_out({mx1_f1_out}), .func2_out({mx1_f2_out}), .func3_out({mx1_f3_out}), 
            .func0_dir({mx1_f0_dir}), .func1_dir({mx1_f1_dir}), .func2_dir({mx1_f2_dir}), 
            .func3_dir({mx1_f3_dir}), .addr({32'b00000000000000000000000000000100}), 
            .sys_w_addr({sys_w_addr}), .sys_r_addr({sys_r_addr}), .sys_w_line({sys_w_line}), 
            .sys_r_line({sys_r_line}), .sys_w(sys_w), .sys_r(sys_r), .rst(rst), 
            .clk(clk));   // test_periph_assembly.v(64)
    gpio_mux mx2 (.pins({pins[95:64]}), .func0_in({g2_in}), .func0_out({mx2_f0_out}), 
            .func1_out({mx2_f1_out}), .func2_out({mx2_f2_out}), .func3_out({mx2_f3_out}), 
            .func0_dir({mx2_f0_dir}), .func1_dir({mx2_f1_dir}), .func2_dir({mx2_f2_dir}), 
            .func3_dir({mx2_f3_dir}), .addr({32'b00000000000000000000000000000110}), 
            .sys_w_addr({sys_w_addr}), .sys_r_addr({sys_r_addr}), .sys_w_line({sys_w_line}), 
            .sys_r_line({sys_r_line}), .sys_w(sys_w), .sys_r(sys_r), .rst(rst), 
            .clk(clk));   // test_periph_assembly.v(65)
    gpio_mux mx3 (.pins({pins[127:96]}), .func0_in({g3_in}), .func0_out({mx3_f0_out}), 
            .func1_out({mx3_f1_out}), .func2_out({mx3_f2_out}), .func3_out({mx3_f3_out}), 
            .func0_dir({mx3_f0_dir}), .func1_dir({mx3_f1_dir}), .func2_dir({mx3_f2_dir}), 
            .func3_dir({mx3_f3_dir}), .addr({32'b00000000000000000000000000001000}), 
            .sys_w_addr({sys_w_addr}), .sys_r_addr({sys_r_addr}), .sys_w_line({sys_w_line}), 
            .sys_r_line({sys_r_line}), .sys_w(sys_w), .sys_r(sys_r), .rst(rst), 
            .clk(clk));   // test_periph_assembly.v(66)
    
endmodule

//
// Verific Verilog Description of module gpio
//

module gpio (gpio_out, gpio_in, gpio_dir, addr, sys_w_addr, sys_r_addr, 
            sys_w_line, sys_r_line, sys_w, sys_r, rst, clk);   // gpio.v(3)
    output [31:0]gpio_out;   // gpio.v(6)
    input [31:0]gpio_in;   // gpio.v(5)
    output [31:0]gpio_dir;   // gpio.v(7)
    input [31:0]addr;   // gpio.v(10)
    input [31:0]sys_w_addr;   // gpio.v(13)
    input [31:0]sys_r_addr;   // gpio.v(14)
    input [31:0]sys_w_line;   // gpio.v(15)
    output [31:0]sys_r_line;   // gpio.v(16)
    input sys_w;   // gpio.v(17)
    input sys_r;   // gpio.v(18)
    input rst;   // gpio.v(22)
    input clk;   // gpio.v(21)
    
    
    wire n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
        n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, 
        n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, 
        n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
        n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, 
        n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, 
        n66, n67, n68, n133, n134, n135, n136, n137, n138, 
        n139, n140, n141, n142, n143, n144, n145, n146, n147, 
        n148, n149, n150, n151, n152, n153, n154, n155, n156, 
        n157, n158, n159, n160, n161, n162, n163, n164, n165, 
        n166, n167, n168, n169, n170, n171, n172, n173, n174, 
        n175, n176, n177, n178, n179, n180, n181, n182, n183, 
        n184, n185, n186, n187, n188, n189, n190, n191, n192, 
        n193, n194, n195, n196, n197, n198, n199, n200, n201, 
        n202, n203, n204, n205, n206, n207, n208, n209, n210, 
        n211, n212, n213, n214, n215, n216, n217, n218, n219, 
        n220, n221, n222, n223, n224, n225, n226, n227, n228, 
        n229, n230, n231, n232, n233, n234, n235, n236, n237, 
        n238, n239, n240, n241, n242, n243, n244, n245, n246, 
        n247, n248, n249, n250, n251, n252, n253, n254, n255, 
        n256, n257, n258, n259, n260, n261, n262, n263, n264, 
        n265, n266, n267, n268, n269, n270, n271, n272, n273, 
        n274, n275, n276, n277, n278, n279, n280, n281, n282, 
        n283, n284, n285, n286, n287, n288, n289, n290, n291, 
        n292, n293, n294, n295, n296, n297, n298, n299, n300, 
        n301, n302, n303, n304, n305, n306, n307, n308, n309, 
        n310, n311, n312, n313, n314, n315, n316, n317, n318, 
        n319, n320, n321, n322, n323, n324, n325, n326, n327, 
        n328, n329, n330, n331, n332, n333, n334, n335, n336, 
        n337, n338, n339, n340, n341, n342, n343, n344, n345, 
        n346, n347, n348, n349, n350, n351, n352, n353, n354, 
        n355, n356, n421, n422, n423, n424, n425, n426, n427, 
        n428, n429, n430, n431, n432, n433, n434, n435, n436, 
        n437, n438, n439, n440, n441, n442, n443, n444, n445, 
        n446, n447, n448, n449, n450, n451, n452, n457, n739;
    
    xor (n5, sys_r_addr[1], addr[1]) ;   // gpio.v(40)
    xor (n6, sys_r_addr[2], addr[2]) ;   // gpio.v(40)
    xor (n7, sys_r_addr[3], addr[3]) ;   // gpio.v(40)
    xor (n8, sys_r_addr[4], addr[4]) ;   // gpio.v(40)
    xor (n9, sys_r_addr[5], addr[5]) ;   // gpio.v(40)
    xor (n10, sys_r_addr[6], addr[6]) ;   // gpio.v(40)
    xor (n11, sys_r_addr[7], addr[7]) ;   // gpio.v(40)
    xor (n12, sys_r_addr[8], addr[8]) ;   // gpio.v(40)
    xor (n13, sys_r_addr[9], addr[9]) ;   // gpio.v(40)
    xor (n14, sys_r_addr[10], addr[10]) ;   // gpio.v(40)
    xor (n15, sys_r_addr[11], addr[11]) ;   // gpio.v(40)
    xor (n16, sys_r_addr[12], addr[12]) ;   // gpio.v(40)
    xor (n17, sys_r_addr[13], addr[13]) ;   // gpio.v(40)
    xor (n18, sys_r_addr[14], addr[14]) ;   // gpio.v(40)
    xor (n19, sys_r_addr[15], addr[15]) ;   // gpio.v(40)
    xor (n20, sys_r_addr[16], addr[16]) ;   // gpio.v(40)
    xor (n21, sys_r_addr[17], addr[17]) ;   // gpio.v(40)
    xor (n22, sys_r_addr[18], addr[18]) ;   // gpio.v(40)
    xor (n23, sys_r_addr[19], addr[19]) ;   // gpio.v(40)
    xor (n24, sys_r_addr[20], addr[20]) ;   // gpio.v(40)
    xor (n25, sys_r_addr[21], addr[21]) ;   // gpio.v(40)
    xor (n26, sys_r_addr[22], addr[22]) ;   // gpio.v(40)
    xor (n27, sys_r_addr[23], addr[23]) ;   // gpio.v(40)
    xor (n28, sys_r_addr[24], addr[24]) ;   // gpio.v(40)
    xor (n29, sys_r_addr[25], addr[25]) ;   // gpio.v(40)
    xor (n30, sys_r_addr[26], addr[26]) ;   // gpio.v(40)
    xor (n31, sys_r_addr[27], addr[27]) ;   // gpio.v(40)
    xor (n32, sys_r_addr[28], addr[28]) ;   // gpio.v(40)
    xor (n33, sys_r_addr[29], addr[29]) ;   // gpio.v(40)
    xor (n34, sys_r_addr[30], addr[30]) ;   // gpio.v(40)
    xor (n35, sys_r_addr[31], addr[31]) ;   // gpio.v(40)
    nor (n36, n35, n34, n33, n32, n31, n30, n29, n28, n27, 
        n26, n25, n24, n23, n22, n21, n20, n19, n18, n17, 
        n16, n15, n14, n13, n12, n11, n10, n9, n8, n7, n6, 
        n5) ;   // gpio.v(40)
    assign n37 = sys_r_addr[0] ? gpio_dir[31] : gpio_in[31];   // gpio.v(43)
    assign n38 = sys_r_addr[0] ? gpio_dir[30] : gpio_in[30];   // gpio.v(43)
    assign n39 = sys_r_addr[0] ? gpio_dir[29] : gpio_in[29];   // gpio.v(43)
    assign n40 = sys_r_addr[0] ? gpio_dir[28] : gpio_in[28];   // gpio.v(43)
    assign n41 = sys_r_addr[0] ? gpio_dir[27] : gpio_in[27];   // gpio.v(43)
    assign n42 = sys_r_addr[0] ? gpio_dir[26] : gpio_in[26];   // gpio.v(43)
    assign n43 = sys_r_addr[0] ? gpio_dir[25] : gpio_in[25];   // gpio.v(43)
    assign n44 = sys_r_addr[0] ? gpio_dir[24] : gpio_in[24];   // gpio.v(43)
    assign n45 = sys_r_addr[0] ? gpio_dir[23] : gpio_in[23];   // gpio.v(43)
    assign n46 = sys_r_addr[0] ? gpio_dir[22] : gpio_in[22];   // gpio.v(43)
    assign n47 = sys_r_addr[0] ? gpio_dir[21] : gpio_in[21];   // gpio.v(43)
    assign n48 = sys_r_addr[0] ? gpio_dir[20] : gpio_in[20];   // gpio.v(43)
    assign n49 = sys_r_addr[0] ? gpio_dir[19] : gpio_in[19];   // gpio.v(43)
    assign n50 = sys_r_addr[0] ? gpio_dir[18] : gpio_in[18];   // gpio.v(43)
    assign n51 = sys_r_addr[0] ? gpio_dir[17] : gpio_in[17];   // gpio.v(43)
    assign n52 = sys_r_addr[0] ? gpio_dir[16] : gpio_in[16];   // gpio.v(43)
    assign n53 = sys_r_addr[0] ? gpio_dir[15] : gpio_in[15];   // gpio.v(43)
    assign n54 = sys_r_addr[0] ? gpio_dir[14] : gpio_in[14];   // gpio.v(43)
    assign n55 = sys_r_addr[0] ? gpio_dir[13] : gpio_in[13];   // gpio.v(43)
    assign n56 = sys_r_addr[0] ? gpio_dir[12] : gpio_in[12];   // gpio.v(43)
    assign n57 = sys_r_addr[0] ? gpio_dir[11] : gpio_in[11];   // gpio.v(43)
    assign n58 = sys_r_addr[0] ? gpio_dir[10] : gpio_in[10];   // gpio.v(43)
    assign n59 = sys_r_addr[0] ? gpio_dir[9] : gpio_in[9];   // gpio.v(43)
    assign n60 = sys_r_addr[0] ? gpio_dir[8] : gpio_in[8];   // gpio.v(43)
    assign n61 = sys_r_addr[0] ? gpio_dir[7] : gpio_in[7];   // gpio.v(43)
    assign n62 = sys_r_addr[0] ? gpio_dir[6] : gpio_in[6];   // gpio.v(43)
    assign n63 = sys_r_addr[0] ? gpio_dir[5] : gpio_in[5];   // gpio.v(43)
    assign n64 = sys_r_addr[0] ? gpio_dir[4] : gpio_in[4];   // gpio.v(43)
    assign n65 = sys_r_addr[0] ? gpio_dir[3] : gpio_in[3];   // gpio.v(43)
    assign n66 = sys_r_addr[0] ? gpio_dir[2] : gpio_in[2];   // gpio.v(43)
    assign n67 = sys_r_addr[0] ? gpio_dir[1] : gpio_in[1];   // gpio.v(43)
    assign n68 = sys_r_addr[0] ? gpio_dir[0] : gpio_in[0];   // gpio.v(43)
    xor (n133, sys_w_addr[1], addr[1]) ;   // gpio.v(53)
    xor (n134, sys_w_addr[2], addr[2]) ;   // gpio.v(53)
    xor (n135, sys_w_addr[3], addr[3]) ;   // gpio.v(53)
    xor (n136, sys_w_addr[4], addr[4]) ;   // gpio.v(53)
    xor (n137, sys_w_addr[5], addr[5]) ;   // gpio.v(53)
    xor (n138, sys_w_addr[6], addr[6]) ;   // gpio.v(53)
    xor (n139, sys_w_addr[7], addr[7]) ;   // gpio.v(53)
    xor (n140, sys_w_addr[8], addr[8]) ;   // gpio.v(53)
    xor (n141, sys_w_addr[9], addr[9]) ;   // gpio.v(53)
    xor (n142, sys_w_addr[10], addr[10]) ;   // gpio.v(53)
    xor (n143, sys_w_addr[11], addr[11]) ;   // gpio.v(53)
    xor (n144, sys_w_addr[12], addr[12]) ;   // gpio.v(53)
    xor (n145, sys_w_addr[13], addr[13]) ;   // gpio.v(53)
    xor (n146, sys_w_addr[14], addr[14]) ;   // gpio.v(53)
    xor (n147, sys_w_addr[15], addr[15]) ;   // gpio.v(53)
    xor (n148, sys_w_addr[16], addr[16]) ;   // gpio.v(53)
    xor (n149, sys_w_addr[17], addr[17]) ;   // gpio.v(53)
    xor (n150, sys_w_addr[18], addr[18]) ;   // gpio.v(53)
    xor (n151, sys_w_addr[19], addr[19]) ;   // gpio.v(53)
    xor (n152, sys_w_addr[20], addr[20]) ;   // gpio.v(53)
    xor (n153, sys_w_addr[21], addr[21]) ;   // gpio.v(53)
    xor (n154, sys_w_addr[22], addr[22]) ;   // gpio.v(53)
    xor (n155, sys_w_addr[23], addr[23]) ;   // gpio.v(53)
    xor (n156, sys_w_addr[24], addr[24]) ;   // gpio.v(53)
    xor (n157, sys_w_addr[25], addr[25]) ;   // gpio.v(53)
    xor (n158, sys_w_addr[26], addr[26]) ;   // gpio.v(53)
    xor (n159, sys_w_addr[27], addr[27]) ;   // gpio.v(53)
    xor (n160, sys_w_addr[28], addr[28]) ;   // gpio.v(53)
    xor (n161, sys_w_addr[29], addr[29]) ;   // gpio.v(53)
    xor (n162, sys_w_addr[30], addr[30]) ;   // gpio.v(53)
    xor (n163, sys_w_addr[31], addr[31]) ;   // gpio.v(53)
    nor (n164, n163, n162, n161, n160, n159, n158, n157, n156, 
        n155, n154, n153, n152, n151, n150, n149, n148, n147, 
        n146, n145, n144, n143, n142, n141, n140, n139, n138, 
        n137, n136, n135, n134, n133) ;   // gpio.v(53)
    assign n165 = sys_w_addr[0] ? sys_w_line[31] : gpio_dir[31];   // gpio.v(56)
    assign n166 = sys_w_addr[0] ? sys_w_line[30] : gpio_dir[30];   // gpio.v(56)
    assign n167 = sys_w_addr[0] ? sys_w_line[29] : gpio_dir[29];   // gpio.v(56)
    assign n168 = sys_w_addr[0] ? sys_w_line[28] : gpio_dir[28];   // gpio.v(56)
    assign n169 = sys_w_addr[0] ? sys_w_line[27] : gpio_dir[27];   // gpio.v(56)
    assign n170 = sys_w_addr[0] ? sys_w_line[26] : gpio_dir[26];   // gpio.v(56)
    assign n171 = sys_w_addr[0] ? sys_w_line[25] : gpio_dir[25];   // gpio.v(56)
    assign n172 = sys_w_addr[0] ? sys_w_line[24] : gpio_dir[24];   // gpio.v(56)
    assign n173 = sys_w_addr[0] ? sys_w_line[23] : gpio_dir[23];   // gpio.v(56)
    assign n174 = sys_w_addr[0] ? sys_w_line[22] : gpio_dir[22];   // gpio.v(56)
    assign n175 = sys_w_addr[0] ? sys_w_line[21] : gpio_dir[21];   // gpio.v(56)
    assign n176 = sys_w_addr[0] ? sys_w_line[20] : gpio_dir[20];   // gpio.v(56)
    assign n177 = sys_w_addr[0] ? sys_w_line[19] : gpio_dir[19];   // gpio.v(56)
    assign n178 = sys_w_addr[0] ? sys_w_line[18] : gpio_dir[18];   // gpio.v(56)
    assign n179 = sys_w_addr[0] ? sys_w_line[17] : gpio_dir[17];   // gpio.v(56)
    assign n180 = sys_w_addr[0] ? sys_w_line[16] : gpio_dir[16];   // gpio.v(56)
    assign n181 = sys_w_addr[0] ? sys_w_line[15] : gpio_dir[15];   // gpio.v(56)
    assign n182 = sys_w_addr[0] ? sys_w_line[14] : gpio_dir[14];   // gpio.v(56)
    assign n183 = sys_w_addr[0] ? sys_w_line[13] : gpio_dir[13];   // gpio.v(56)
    assign n184 = sys_w_addr[0] ? sys_w_line[12] : gpio_dir[12];   // gpio.v(56)
    assign n185 = sys_w_addr[0] ? sys_w_line[11] : gpio_dir[11];   // gpio.v(56)
    assign n186 = sys_w_addr[0] ? sys_w_line[10] : gpio_dir[10];   // gpio.v(56)
    assign n187 = sys_w_addr[0] ? sys_w_line[9] : gpio_dir[9];   // gpio.v(56)
    assign n188 = sys_w_addr[0] ? sys_w_line[8] : gpio_dir[8];   // gpio.v(56)
    assign n189 = sys_w_addr[0] ? sys_w_line[7] : gpio_dir[7];   // gpio.v(56)
    assign n190 = sys_w_addr[0] ? sys_w_line[6] : gpio_dir[6];   // gpio.v(56)
    assign n191 = sys_w_addr[0] ? sys_w_line[5] : gpio_dir[5];   // gpio.v(56)
    assign n192 = sys_w_addr[0] ? sys_w_line[4] : gpio_dir[4];   // gpio.v(56)
    assign n193 = sys_w_addr[0] ? sys_w_line[3] : gpio_dir[3];   // gpio.v(56)
    assign n194 = sys_w_addr[0] ? sys_w_line[2] : gpio_dir[2];   // gpio.v(56)
    assign n195 = sys_w_addr[0] ? sys_w_line[1] : gpio_dir[1];   // gpio.v(56)
    assign n196 = sys_w_addr[0] ? sys_w_line[0] : gpio_dir[0];   // gpio.v(56)
    assign n197 = sys_w_addr[0] ? gpio_out[31] : sys_w_line[31];   // gpio.v(56)
    assign n198 = sys_w_addr[0] ? gpio_out[30] : sys_w_line[30];   // gpio.v(56)
    assign n199 = sys_w_addr[0] ? gpio_out[29] : sys_w_line[29];   // gpio.v(56)
    assign n200 = sys_w_addr[0] ? gpio_out[28] : sys_w_line[28];   // gpio.v(56)
    assign n201 = sys_w_addr[0] ? gpio_out[27] : sys_w_line[27];   // gpio.v(56)
    assign n202 = sys_w_addr[0] ? gpio_out[26] : sys_w_line[26];   // gpio.v(56)
    assign n203 = sys_w_addr[0] ? gpio_out[25] : sys_w_line[25];   // gpio.v(56)
    assign n204 = sys_w_addr[0] ? gpio_out[24] : sys_w_line[24];   // gpio.v(56)
    assign n205 = sys_w_addr[0] ? gpio_out[23] : sys_w_line[23];   // gpio.v(56)
    assign n206 = sys_w_addr[0] ? gpio_out[22] : sys_w_line[22];   // gpio.v(56)
    assign n207 = sys_w_addr[0] ? gpio_out[21] : sys_w_line[21];   // gpio.v(56)
    assign n208 = sys_w_addr[0] ? gpio_out[20] : sys_w_line[20];   // gpio.v(56)
    assign n209 = sys_w_addr[0] ? gpio_out[19] : sys_w_line[19];   // gpio.v(56)
    assign n210 = sys_w_addr[0] ? gpio_out[18] : sys_w_line[18];   // gpio.v(56)
    assign n211 = sys_w_addr[0] ? gpio_out[17] : sys_w_line[17];   // gpio.v(56)
    assign n212 = sys_w_addr[0] ? gpio_out[16] : sys_w_line[16];   // gpio.v(56)
    assign n213 = sys_w_addr[0] ? gpio_out[15] : sys_w_line[15];   // gpio.v(56)
    assign n214 = sys_w_addr[0] ? gpio_out[14] : sys_w_line[14];   // gpio.v(56)
    assign n215 = sys_w_addr[0] ? gpio_out[13] : sys_w_line[13];   // gpio.v(56)
    assign n216 = sys_w_addr[0] ? gpio_out[12] : sys_w_line[12];   // gpio.v(56)
    assign n217 = sys_w_addr[0] ? gpio_out[11] : sys_w_line[11];   // gpio.v(56)
    assign n218 = sys_w_addr[0] ? gpio_out[10] : sys_w_line[10];   // gpio.v(56)
    assign n219 = sys_w_addr[0] ? gpio_out[9] : sys_w_line[9];   // gpio.v(56)
    assign n220 = sys_w_addr[0] ? gpio_out[8] : sys_w_line[8];   // gpio.v(56)
    assign n221 = sys_w_addr[0] ? gpio_out[7] : sys_w_line[7];   // gpio.v(56)
    assign n222 = sys_w_addr[0] ? gpio_out[6] : sys_w_line[6];   // gpio.v(56)
    assign n223 = sys_w_addr[0] ? gpio_out[5] : sys_w_line[5];   // gpio.v(56)
    assign n224 = sys_w_addr[0] ? gpio_out[4] : sys_w_line[4];   // gpio.v(56)
    assign n225 = sys_w_addr[0] ? gpio_out[3] : sys_w_line[3];   // gpio.v(56)
    assign n226 = sys_w_addr[0] ? gpio_out[2] : sys_w_line[2];   // gpio.v(56)
    assign n227 = sys_w_addr[0] ? gpio_out[1] : sys_w_line[1];   // gpio.v(56)
    assign n228 = sys_w_addr[0] ? gpio_out[0] : sys_w_line[0];   // gpio.v(56)
    assign n229 = n164 ? n165 : gpio_dir[31];   // gpio.v(53)
    assign n230 = n164 ? n166 : gpio_dir[30];   // gpio.v(53)
    assign n231 = n164 ? n167 : gpio_dir[29];   // gpio.v(53)
    assign n232 = n164 ? n168 : gpio_dir[28];   // gpio.v(53)
    assign n233 = n164 ? n169 : gpio_dir[27];   // gpio.v(53)
    assign n234 = n164 ? n170 : gpio_dir[26];   // gpio.v(53)
    assign n235 = n164 ? n171 : gpio_dir[25];   // gpio.v(53)
    assign n236 = n164 ? n172 : gpio_dir[24];   // gpio.v(53)
    assign n237 = n164 ? n173 : gpio_dir[23];   // gpio.v(53)
    assign n238 = n164 ? n174 : gpio_dir[22];   // gpio.v(53)
    assign n239 = n164 ? n175 : gpio_dir[21];   // gpio.v(53)
    assign n240 = n164 ? n176 : gpio_dir[20];   // gpio.v(53)
    assign n241 = n164 ? n177 : gpio_dir[19];   // gpio.v(53)
    assign n242 = n164 ? n178 : gpio_dir[18];   // gpio.v(53)
    assign n243 = n164 ? n179 : gpio_dir[17];   // gpio.v(53)
    assign n244 = n164 ? n180 : gpio_dir[16];   // gpio.v(53)
    assign n245 = n164 ? n181 : gpio_dir[15];   // gpio.v(53)
    assign n246 = n164 ? n182 : gpio_dir[14];   // gpio.v(53)
    assign n247 = n164 ? n183 : gpio_dir[13];   // gpio.v(53)
    assign n248 = n164 ? n184 : gpio_dir[12];   // gpio.v(53)
    assign n249 = n164 ? n185 : gpio_dir[11];   // gpio.v(53)
    assign n250 = n164 ? n186 : gpio_dir[10];   // gpio.v(53)
    assign n251 = n164 ? n187 : gpio_dir[9];   // gpio.v(53)
    assign n252 = n164 ? n188 : gpio_dir[8];   // gpio.v(53)
    assign n253 = n164 ? n189 : gpio_dir[7];   // gpio.v(53)
    assign n254 = n164 ? n190 : gpio_dir[6];   // gpio.v(53)
    assign n255 = n164 ? n191 : gpio_dir[5];   // gpio.v(53)
    assign n256 = n164 ? n192 : gpio_dir[4];   // gpio.v(53)
    assign n257 = n164 ? n193 : gpio_dir[3];   // gpio.v(53)
    assign n258 = n164 ? n194 : gpio_dir[2];   // gpio.v(53)
    assign n259 = n164 ? n195 : gpio_dir[1];   // gpio.v(53)
    assign n260 = n164 ? n196 : gpio_dir[0];   // gpio.v(53)
    assign n261 = n164 ? n197 : gpio_out[31];   // gpio.v(53)
    assign n262 = n164 ? n198 : gpio_out[30];   // gpio.v(53)
    assign n263 = n164 ? n199 : gpio_out[29];   // gpio.v(53)
    assign n264 = n164 ? n200 : gpio_out[28];   // gpio.v(53)
    assign n265 = n164 ? n201 : gpio_out[27];   // gpio.v(53)
    assign n266 = n164 ? n202 : gpio_out[26];   // gpio.v(53)
    assign n267 = n164 ? n203 : gpio_out[25];   // gpio.v(53)
    assign n268 = n164 ? n204 : gpio_out[24];   // gpio.v(53)
    assign n269 = n164 ? n205 : gpio_out[23];   // gpio.v(53)
    assign n270 = n164 ? n206 : gpio_out[22];   // gpio.v(53)
    assign n271 = n164 ? n207 : gpio_out[21];   // gpio.v(53)
    assign n272 = n164 ? n208 : gpio_out[20];   // gpio.v(53)
    assign n273 = n164 ? n209 : gpio_out[19];   // gpio.v(53)
    assign n274 = n164 ? n210 : gpio_out[18];   // gpio.v(53)
    assign n275 = n164 ? n211 : gpio_out[17];   // gpio.v(53)
    assign n276 = n164 ? n212 : gpio_out[16];   // gpio.v(53)
    assign n277 = n164 ? n213 : gpio_out[15];   // gpio.v(53)
    assign n278 = n164 ? n214 : gpio_out[14];   // gpio.v(53)
    assign n279 = n164 ? n215 : gpio_out[13];   // gpio.v(53)
    assign n280 = n164 ? n216 : gpio_out[12];   // gpio.v(53)
    assign n281 = n164 ? n217 : gpio_out[11];   // gpio.v(53)
    assign n282 = n164 ? n218 : gpio_out[10];   // gpio.v(53)
    assign n283 = n164 ? n219 : gpio_out[9];   // gpio.v(53)
    assign n284 = n164 ? n220 : gpio_out[8];   // gpio.v(53)
    assign n285 = n164 ? n221 : gpio_out[7];   // gpio.v(53)
    assign n286 = n164 ? n222 : gpio_out[6];   // gpio.v(53)
    assign n287 = n164 ? n223 : gpio_out[5];   // gpio.v(53)
    assign n288 = n164 ? n224 : gpio_out[4];   // gpio.v(53)
    assign n289 = n164 ? n225 : gpio_out[3];   // gpio.v(53)
    assign n290 = n164 ? n226 : gpio_out[2];   // gpio.v(53)
    assign n291 = n164 ? n227 : gpio_out[1];   // gpio.v(53)
    assign n292 = n164 ? n228 : gpio_out[0];   // gpio.v(53)
    assign n293 = sys_w ? n229 : gpio_dir[31];   // gpio.v(52)
    assign n294 = sys_w ? n230 : gpio_dir[30];   // gpio.v(52)
    assign n295 = sys_w ? n231 : gpio_dir[29];   // gpio.v(52)
    assign n296 = sys_w ? n232 : gpio_dir[28];   // gpio.v(52)
    assign n297 = sys_w ? n233 : gpio_dir[27];   // gpio.v(52)
    assign n298 = sys_w ? n234 : gpio_dir[26];   // gpio.v(52)
    assign n299 = sys_w ? n235 : gpio_dir[25];   // gpio.v(52)
    assign n300 = sys_w ? n236 : gpio_dir[24];   // gpio.v(52)
    assign n301 = sys_w ? n237 : gpio_dir[23];   // gpio.v(52)
    assign n302 = sys_w ? n238 : gpio_dir[22];   // gpio.v(52)
    assign n303 = sys_w ? n239 : gpio_dir[21];   // gpio.v(52)
    assign n304 = sys_w ? n240 : gpio_dir[20];   // gpio.v(52)
    assign n305 = sys_w ? n241 : gpio_dir[19];   // gpio.v(52)
    assign n306 = sys_w ? n242 : gpio_dir[18];   // gpio.v(52)
    assign n307 = sys_w ? n243 : gpio_dir[17];   // gpio.v(52)
    assign n308 = sys_w ? n244 : gpio_dir[16];   // gpio.v(52)
    assign n309 = sys_w ? n245 : gpio_dir[15];   // gpio.v(52)
    assign n310 = sys_w ? n246 : gpio_dir[14];   // gpio.v(52)
    assign n311 = sys_w ? n247 : gpio_dir[13];   // gpio.v(52)
    assign n312 = sys_w ? n248 : gpio_dir[12];   // gpio.v(52)
    assign n313 = sys_w ? n249 : gpio_dir[11];   // gpio.v(52)
    assign n314 = sys_w ? n250 : gpio_dir[10];   // gpio.v(52)
    assign n315 = sys_w ? n251 : gpio_dir[9];   // gpio.v(52)
    assign n316 = sys_w ? n252 : gpio_dir[8];   // gpio.v(52)
    assign n317 = sys_w ? n253 : gpio_dir[7];   // gpio.v(52)
    assign n318 = sys_w ? n254 : gpio_dir[6];   // gpio.v(52)
    assign n319 = sys_w ? n255 : gpio_dir[5];   // gpio.v(52)
    assign n320 = sys_w ? n256 : gpio_dir[4];   // gpio.v(52)
    assign n321 = sys_w ? n257 : gpio_dir[3];   // gpio.v(52)
    assign n322 = sys_w ? n258 : gpio_dir[2];   // gpio.v(52)
    assign n323 = sys_w ? n259 : gpio_dir[1];   // gpio.v(52)
    assign n324 = sys_w ? n260 : gpio_dir[0];   // gpio.v(52)
    assign n325 = sys_w ? n261 : gpio_out[31];   // gpio.v(52)
    assign n326 = sys_w ? n262 : gpio_out[30];   // gpio.v(52)
    assign n327 = sys_w ? n263 : gpio_out[29];   // gpio.v(52)
    assign n328 = sys_w ? n264 : gpio_out[28];   // gpio.v(52)
    assign n329 = sys_w ? n265 : gpio_out[27];   // gpio.v(52)
    assign n330 = sys_w ? n266 : gpio_out[26];   // gpio.v(52)
    assign n331 = sys_w ? n267 : gpio_out[25];   // gpio.v(52)
    assign n332 = sys_w ? n268 : gpio_out[24];   // gpio.v(52)
    assign n333 = sys_w ? n269 : gpio_out[23];   // gpio.v(52)
    assign n334 = sys_w ? n270 : gpio_out[22];   // gpio.v(52)
    assign n335 = sys_w ? n271 : gpio_out[21];   // gpio.v(52)
    assign n336 = sys_w ? n272 : gpio_out[20];   // gpio.v(52)
    assign n337 = sys_w ? n273 : gpio_out[19];   // gpio.v(52)
    assign n338 = sys_w ? n274 : gpio_out[18];   // gpio.v(52)
    assign n339 = sys_w ? n275 : gpio_out[17];   // gpio.v(52)
    assign n340 = sys_w ? n276 : gpio_out[16];   // gpio.v(52)
    assign n341 = sys_w ? n277 : gpio_out[15];   // gpio.v(52)
    assign n342 = sys_w ? n278 : gpio_out[14];   // gpio.v(52)
    assign n343 = sys_w ? n279 : gpio_out[13];   // gpio.v(52)
    assign n344 = sys_w ? n280 : gpio_out[12];   // gpio.v(52)
    assign n345 = sys_w ? n281 : gpio_out[11];   // gpio.v(52)
    assign n346 = sys_w ? n282 : gpio_out[10];   // gpio.v(52)
    assign n347 = sys_w ? n283 : gpio_out[9];   // gpio.v(52)
    assign n348 = sys_w ? n284 : gpio_out[8];   // gpio.v(52)
    assign n349 = sys_w ? n285 : gpio_out[7];   // gpio.v(52)
    assign n350 = sys_w ? n286 : gpio_out[6];   // gpio.v(52)
    assign n351 = sys_w ? n287 : gpio_out[5];   // gpio.v(52)
    assign n352 = sys_w ? n288 : gpio_out[4];   // gpio.v(52)
    assign n353 = sys_w ? n289 : gpio_out[3];   // gpio.v(52)
    assign n354 = sys_w ? n290 : gpio_out[2];   // gpio.v(52)
    assign n355 = sys_w ? n291 : gpio_out[1];   // gpio.v(52)
    assign n356 = sys_w ? n292 : gpio_out[0];   // gpio.v(52)
    VERIFIC_DFFRS i358 (.d(n294), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[30]));   // gpio.v(37)
    VERIFIC_DFFRS i359 (.d(n295), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[29]));   // gpio.v(37)
    VERIFIC_DFFRS i360 (.d(n296), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[28]));   // gpio.v(37)
    VERIFIC_DFFRS i361 (.d(n297), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[27]));   // gpio.v(37)
    VERIFIC_DFFRS i362 (.d(n298), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[26]));   // gpio.v(37)
    VERIFIC_DFFRS i363 (.d(n299), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[25]));   // gpio.v(37)
    VERIFIC_DFFRS i364 (.d(n300), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[24]));   // gpio.v(37)
    VERIFIC_DFFRS i365 (.d(n301), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[23]));   // gpio.v(37)
    VERIFIC_DFFRS i366 (.d(n302), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[22]));   // gpio.v(37)
    VERIFIC_DFFRS i367 (.d(n303), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[21]));   // gpio.v(37)
    VERIFIC_DFFRS i368 (.d(n304), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[20]));   // gpio.v(37)
    VERIFIC_DFFRS i369 (.d(n305), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[19]));   // gpio.v(37)
    VERIFIC_DFFRS i370 (.d(n306), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[18]));   // gpio.v(37)
    VERIFIC_DFFRS i371 (.d(n307), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[17]));   // gpio.v(37)
    VERIFIC_DFFRS i372 (.d(n308), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[16]));   // gpio.v(37)
    VERIFIC_DFFRS i373 (.d(n309), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[15]));   // gpio.v(37)
    VERIFIC_DFFRS i374 (.d(n310), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[14]));   // gpio.v(37)
    VERIFIC_DFFRS i375 (.d(n311), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[13]));   // gpio.v(37)
    VERIFIC_DFFRS i376 (.d(n312), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[12]));   // gpio.v(37)
    VERIFIC_DFFRS i377 (.d(n313), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[11]));   // gpio.v(37)
    VERIFIC_DFFRS i378 (.d(n314), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[10]));   // gpio.v(37)
    VERIFIC_DFFRS i379 (.d(n315), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[9]));   // gpio.v(37)
    VERIFIC_DFFRS i380 (.d(n316), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[8]));   // gpio.v(37)
    VERIFIC_DFFRS i381 (.d(n317), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[7]));   // gpio.v(37)
    VERIFIC_DFFRS i382 (.d(n318), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[6]));   // gpio.v(37)
    VERIFIC_DFFRS i383 (.d(n319), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[5]));   // gpio.v(37)
    VERIFIC_DFFRS i384 (.d(n320), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[4]));   // gpio.v(37)
    VERIFIC_DFFRS i385 (.d(n321), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[3]));   // gpio.v(37)
    VERIFIC_DFFRS i386 (.d(n322), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[2]));   // gpio.v(37)
    VERIFIC_DFFRS i387 (.d(n323), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[1]));   // gpio.v(37)
    VERIFIC_DFFRS i388 (.d(n324), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[0]));   // gpio.v(37)
    VERIFIC_DFFRS i389 (.d(n325), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[31]));   // gpio.v(37)
    VERIFIC_DFFRS i390 (.d(n326), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[30]));   // gpio.v(37)
    VERIFIC_DFFRS i391 (.d(n327), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[29]));   // gpio.v(37)
    VERIFIC_DFFRS i392 (.d(n328), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[28]));   // gpio.v(37)
    VERIFIC_DFFRS i393 (.d(n329), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[27]));   // gpio.v(37)
    VERIFIC_DFFRS i394 (.d(n330), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[26]));   // gpio.v(37)
    VERIFIC_DFFRS i395 (.d(n331), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[25]));   // gpio.v(37)
    VERIFIC_DFFRS i396 (.d(n332), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[24]));   // gpio.v(37)
    VERIFIC_DFFRS i397 (.d(n333), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[23]));   // gpio.v(37)
    VERIFIC_DFFRS i398 (.d(n334), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[22]));   // gpio.v(37)
    VERIFIC_DFFRS i399 (.d(n335), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[21]));   // gpio.v(37)
    VERIFIC_DFFRS i400 (.d(n336), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[20]));   // gpio.v(37)
    VERIFIC_DFFRS i401 (.d(n337), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[19]));   // gpio.v(37)
    VERIFIC_DFFRS i402 (.d(n338), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[18]));   // gpio.v(37)
    VERIFIC_DFFRS i403 (.d(n339), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[17]));   // gpio.v(37)
    VERIFIC_DFFRS i404 (.d(n340), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[16]));   // gpio.v(37)
    VERIFIC_DFFRS i405 (.d(n341), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[15]));   // gpio.v(37)
    VERIFIC_DFFRS i406 (.d(n342), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[14]));   // gpio.v(37)
    VERIFIC_DFFRS i407 (.d(n343), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[13]));   // gpio.v(37)
    VERIFIC_DFFRS i408 (.d(n344), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[12]));   // gpio.v(37)
    VERIFIC_DFFRS i409 (.d(n345), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[11]));   // gpio.v(37)
    VERIFIC_DFFRS i410 (.d(n346), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[10]));   // gpio.v(37)
    VERIFIC_DFFRS i411 (.d(n347), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[9]));   // gpio.v(37)
    VERIFIC_DFFRS i412 (.d(n348), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[8]));   // gpio.v(37)
    VERIFIC_DFFRS i413 (.d(n349), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[7]));   // gpio.v(37)
    VERIFIC_DFFRS i414 (.d(n350), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[6]));   // gpio.v(37)
    VERIFIC_DFFRS i415 (.d(n351), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[5]));   // gpio.v(37)
    VERIFIC_DFFRS i416 (.d(n352), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[4]));   // gpio.v(37)
    VERIFIC_DFFRS i417 (.d(n353), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[3]));   // gpio.v(37)
    VERIFIC_DFFRS i418 (.d(n354), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[2]));   // gpio.v(37)
    VERIFIC_DFFRS i419 (.d(n355), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[1]));   // gpio.v(37)
    VERIFIC_DFFRS i420 (.d(n356), .clk(clk), .s(1'b0), .r(rst), .q(gpio_out[0]));   // gpio.v(37)
    VERIFIC_DFFRS i422 (.d(n38), .clk(clk), .s(1'b0), .r(rst), .q(n422));   // gpio.v(37)
    VERIFIC_DFFRS i423 (.d(n39), .clk(clk), .s(1'b0), .r(rst), .q(n423));   // gpio.v(37)
    VERIFIC_DFFRS i424 (.d(n40), .clk(clk), .s(1'b0), .r(rst), .q(n424));   // gpio.v(37)
    VERIFIC_DFFRS i425 (.d(n41), .clk(clk), .s(1'b0), .r(rst), .q(n425));   // gpio.v(37)
    VERIFIC_DFFRS i426 (.d(n42), .clk(clk), .s(1'b0), .r(rst), .q(n426));   // gpio.v(37)
    VERIFIC_DFFRS i427 (.d(n43), .clk(clk), .s(1'b0), .r(rst), .q(n427));   // gpio.v(37)
    VERIFIC_DFFRS i428 (.d(n44), .clk(clk), .s(1'b0), .r(rst), .q(n428));   // gpio.v(37)
    VERIFIC_DFFRS i429 (.d(n45), .clk(clk), .s(1'b0), .r(rst), .q(n429));   // gpio.v(37)
    VERIFIC_DFFRS i430 (.d(n46), .clk(clk), .s(1'b0), .r(rst), .q(n430));   // gpio.v(37)
    VERIFIC_DFFRS i431 (.d(n47), .clk(clk), .s(1'b0), .r(rst), .q(n431));   // gpio.v(37)
    VERIFIC_DFFRS i432 (.d(n48), .clk(clk), .s(1'b0), .r(rst), .q(n432));   // gpio.v(37)
    VERIFIC_DFFRS i433 (.d(n49), .clk(clk), .s(1'b0), .r(rst), .q(n433));   // gpio.v(37)
    VERIFIC_DFFRS i434 (.d(n50), .clk(clk), .s(1'b0), .r(rst), .q(n434));   // gpio.v(37)
    VERIFIC_DFFRS i435 (.d(n51), .clk(clk), .s(1'b0), .r(rst), .q(n435));   // gpio.v(37)
    VERIFIC_DFFRS i436 (.d(n52), .clk(clk), .s(1'b0), .r(rst), .q(n436));   // gpio.v(37)
    VERIFIC_DFFRS i437 (.d(n53), .clk(clk), .s(1'b0), .r(rst), .q(n437));   // gpio.v(37)
    VERIFIC_DFFRS i438 (.d(n54), .clk(clk), .s(1'b0), .r(rst), .q(n438));   // gpio.v(37)
    VERIFIC_DFFRS i439 (.d(n55), .clk(clk), .s(1'b0), .r(rst), .q(n439));   // gpio.v(37)
    VERIFIC_DFFRS i440 (.d(n56), .clk(clk), .s(1'b0), .r(rst), .q(n440));   // gpio.v(37)
    VERIFIC_DFFRS i441 (.d(n57), .clk(clk), .s(1'b0), .r(rst), .q(n441));   // gpio.v(37)
    VERIFIC_DFFRS i442 (.d(n58), .clk(clk), .s(1'b0), .r(rst), .q(n442));   // gpio.v(37)
    VERIFIC_DFFRS i443 (.d(n59), .clk(clk), .s(1'b0), .r(rst), .q(n443));   // gpio.v(37)
    VERIFIC_DFFRS i444 (.d(n60), .clk(clk), .s(1'b0), .r(rst), .q(n444));   // gpio.v(37)
    VERIFIC_DFFRS i445 (.d(n61), .clk(clk), .s(1'b0), .r(rst), .q(n445));   // gpio.v(37)
    VERIFIC_DFFRS i446 (.d(n62), .clk(clk), .s(1'b0), .r(rst), .q(n446));   // gpio.v(37)
    VERIFIC_DFFRS i447 (.d(n63), .clk(clk), .s(1'b0), .r(rst), .q(n447));   // gpio.v(37)
    VERIFIC_DFFRS i448 (.d(n64), .clk(clk), .s(1'b0), .r(rst), .q(n448));   // gpio.v(37)
    VERIFIC_DFFRS i449 (.d(n65), .clk(clk), .s(1'b0), .r(rst), .q(n449));   // gpio.v(37)
    VERIFIC_DFFRS i450 (.d(n66), .clk(clk), .s(1'b0), .r(rst), .q(n450));   // gpio.v(37)
    VERIFIC_DFFRS i451 (.d(n67), .clk(clk), .s(1'b0), .r(rst), .q(n451));   // gpio.v(37)
    VERIFIC_DFFRS i452 (.d(n68), .clk(clk), .s(1'b0), .r(rst), .q(n452));   // gpio.v(37)
    and (n457, sys_r, n36) ;   // gpio.v(49)
    assign sys_r_line[31] = n739 ? n421 : 1'bz;   // gpio.v(31)
    assign sys_r_line[30] = n739 ? n422 : 1'bz;   // gpio.v(31)
    assign sys_r_line[29] = n739 ? n423 : 1'bz;   // gpio.v(31)
    assign sys_r_line[28] = n739 ? n424 : 1'bz;   // gpio.v(31)
    assign sys_r_line[27] = n739 ? n425 : 1'bz;   // gpio.v(31)
    assign sys_r_line[26] = n739 ? n426 : 1'bz;   // gpio.v(31)
    assign sys_r_line[25] = n739 ? n427 : 1'bz;   // gpio.v(31)
    assign sys_r_line[24] = n739 ? n428 : 1'bz;   // gpio.v(31)
    assign sys_r_line[23] = n739 ? n429 : 1'bz;   // gpio.v(31)
    assign sys_r_line[22] = n739 ? n430 : 1'bz;   // gpio.v(31)
    assign sys_r_line[21] = n739 ? n431 : 1'bz;   // gpio.v(31)
    assign sys_r_line[20] = n739 ? n432 : 1'bz;   // gpio.v(31)
    assign sys_r_line[19] = n739 ? n433 : 1'bz;   // gpio.v(31)
    assign sys_r_line[18] = n739 ? n434 : 1'bz;   // gpio.v(31)
    assign sys_r_line[17] = n739 ? n435 : 1'bz;   // gpio.v(31)
    assign sys_r_line[16] = n739 ? n436 : 1'bz;   // gpio.v(31)
    assign sys_r_line[15] = n739 ? n437 : 1'bz;   // gpio.v(31)
    assign sys_r_line[14] = n739 ? n438 : 1'bz;   // gpio.v(31)
    assign sys_r_line[13] = n739 ? n439 : 1'bz;   // gpio.v(31)
    assign sys_r_line[12] = n739 ? n440 : 1'bz;   // gpio.v(31)
    assign sys_r_line[11] = n739 ? n441 : 1'bz;   // gpio.v(31)
    assign sys_r_line[10] = n739 ? n442 : 1'bz;   // gpio.v(31)
    assign sys_r_line[9] = n739 ? n443 : 1'bz;   // gpio.v(31)
    assign sys_r_line[8] = n739 ? n444 : 1'bz;   // gpio.v(31)
    assign sys_r_line[7] = n739 ? n445 : 1'bz;   // gpio.v(31)
    assign sys_r_line[6] = n739 ? n446 : 1'bz;   // gpio.v(31)
    assign sys_r_line[5] = n739 ? n447 : 1'bz;   // gpio.v(31)
    assign sys_r_line[4] = n739 ? n448 : 1'bz;   // gpio.v(31)
    assign sys_r_line[3] = n739 ? n449 : 1'bz;   // gpio.v(31)
    assign sys_r_line[2] = n739 ? n450 : 1'bz;   // gpio.v(31)
    VERIFIC_DFFRS i739 (.d(n457), .clk(clk), .s(1'b0), .r(rst), .q(n739));   // gpio.v(37)
    assign sys_r_line[1] = n739 ? n451 : 1'bz;   // gpio.v(31)
    assign sys_r_line[0] = n739 ? n452 : 1'bz;   // gpio.v(31)
    VERIFIC_DFFRS i357 (.d(n293), .clk(clk), .s(1'b0), .r(rst), .q(gpio_dir[31]));   // gpio.v(37)
    VERIFIC_DFFRS i421 (.d(n37), .clk(clk), .s(1'b0), .r(rst), .q(n421));   // gpio.v(37)
    
endmodule

//
// Verific Verilog Description of PRIMITIVE VERIFIC_DFFRS
//

module VERIFIC_DFFRS (d, clk, s, r, q);
    input d;
    input clk;
    input s;
    input r;
    output q;
    reg q ;
    always @(posedge clk or posedge s or posedge r) begin
        if (s) q = 1'b1;
        else if (r) q = 1'b0;
        else q = d;
    end
    
endmodule

//
// Verific Verilog Description of module gpio_mux
//

module gpio_mux (pins, func0_in, func1_in, func2_in, func3_in, func0_out, 
            func1_out, func2_out, func3_out, func0_dir, func1_dir, 
            func2_dir, func3_dir, addr, sys_w_addr, sys_r_addr, sys_w_line, 
            sys_r_line, sys_w, sys_r, rst, clk);   // gpio_mux.v(3)
    inout [31:0]pins;   // gpio_mux.v(4)
    output [31:0]func0_in;   // gpio_mux.v(14)
    output [31:0]func1_in;   // gpio_mux.v(15)
    output [31:0]func2_in;   // gpio_mux.v(16)
    output [31:0]func3_in;   // gpio_mux.v(17)
    input [31:0]func0_out;   // gpio_mux.v(8)
    input [31:0]func1_out;   // gpio_mux.v(9)
    input [31:0]func2_out;   // gpio_mux.v(10)
    input [31:0]func3_out;   // gpio_mux.v(11)
    input [31:0]func0_dir;   // gpio_mux.v(20)
    input [31:0]func1_dir;   // gpio_mux.v(21)
    input [31:0]func2_dir;   // gpio_mux.v(22)
    input [31:0]func3_dir;   // gpio_mux.v(23)
    input [31:0]addr;   // gpio_mux.v(26)
    input [31:0]sys_w_addr;   // gpio_mux.v(29)
    input [31:0]sys_r_addr;   // gpio_mux.v(30)
    input [31:0]sys_w_line;   // gpio_mux.v(31)
    output [31:0]sys_r_line;   // gpio_mux.v(32)
    input sys_w;   // gpio_mux.v(33)
    input sys_r;   // gpio_mux.v(34)
    input rst;   // gpio_mux.v(38)
    input clk;   // gpio_mux.v(37)
    
    wire [1:0]\pin_mux[0].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[0].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[0].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[1].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[1].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[1].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[2].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[2].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[2].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[3].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[3].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[3].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[4].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[4].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[4].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[5].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[5].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[5].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[6].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[6].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[6].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[7].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[7].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[7].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[8].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[8].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[8].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[9].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[9].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[9].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[10].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[10].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[10].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[11].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[11].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[11].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[12].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[12].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[12].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[13].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[13].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[13].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[14].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[14].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[14].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[15].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[15].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[15].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[16].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[16].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[16].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[17].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[17].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[17].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[18].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[18].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[18].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[19].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[19].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[19].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[20].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[20].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[20].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[21].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[21].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[21].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[22].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[22].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[22].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[23].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[23].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[23].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[24].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[24].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[24].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[25].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[25].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[25].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[26].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[26].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[26].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[27].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[27].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[27].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[28].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[28].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[28].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[29].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[29].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[29].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[30].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[30].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[30].pin_dir ;   // gpio_mux.v(49)
    wire [1:0]\pin_mux[31].pin_control ;   // gpio_mux.v(47)
    wire \pin_mux[31].pin_out ;   // gpio_mux.v(48)
    wire \pin_mux[31].pin_dir ;   // gpio_mux.v(49)
    
    wire n4, n5, n6, n7, n8, n9, n10, n17, n18, n33, n34, 
        n35, n36, n37, n38, n39, n46, n47, n62, n63, n64, 
        n65, n66, n67, n68, n75, n76, n91, n92, n93, n94, 
        n95, n96, n97, n104, n105, n120, n121, n122, n123, 
        n124, n125, n126, n133, n134, n149, n150, n151, n152, 
        n153, n154, n155, n162, n163, n178, n179, n180, n181, 
        n182, n183, n184, n191, n192, n207, n208, n209, n210, 
        n211, n212, n213, n220, n221, n236, n237, n238, n239, 
        n240, n241, n242, n249, n250, n265, n266, n267, n268, 
        n269, n270, n271, n278, n279, n294, n295, n296, n297, 
        n298, n299, n300, n307, n308, n323, n324, n325, n326, 
        n327, n328, n329, n336, n337, n352, n353, n354, n355, 
        n356, n357, n358, n365, n366, n381, n382, n383, n384, 
        n385, n386, n387, n394, n395, n410, n411, n412, n413, 
        n414, n415, n416, n423, n424, n439, n440, n441, n442, 
        n443, n444, n445, n452, n453, n468, n469, n470, n471, 
        n472, n473, n474, n481, n482, n497, n498, n499, n500, 
        n501, n502, n503, n510, n511, n526, n527, n528, n529, 
        n530, n531, n532, n539, n540, n555, n556, n557, n558, 
        n559, n560, n561, n568, n569, n584, n585, n586, n587, 
        n588, n589, n590, n597, n598, n613, n614, n615, n616, 
        n617, n618, n619, n626, n627, n642, n643, n644, n645, 
        n646, n647, n648, n655, n656, n671, n672, n673, n674, 
        n675, n676, n677, n684, n685, n700, n701, n702, n703, 
        n704, n705, n706, n713, n714, n729, n730, n731, n732, 
        n733, n734, n735, n742, n743, n758, n759, n760, n761, 
        n762, n763, n764, n771, n772, n787, n788, n789, n790, 
        n791, n792, n793, n800, n801, n816, n817, n818, n819, 
        n820, n821, n822, n829, n830, n845, n846, n847, n848, 
        n849, n850, n851, n858, n859, n874, n875, n876, n877, 
        n878, n879, n880, n887, n888, n903, n904, n905, n906, 
        n907, n908, n909, n916, n917, n933, n934, n935, n936, 
        n937, n938, n939, n940, n941, n942, n943, n944, n945, 
        n946, n947, n948, n949, n950, n951, n952, n953, n954, 
        n955, n956, n957, n958, n959, n960, n961, n962, n963, 
        n964, n965, n966, n967, n968, n969, n970, n971, n972, 
        n973, n974, n975, n976, n977, n978, n979, n980, n981, 
        n982, n983, n984, n985, n986, n987, n988, n989, n990, 
        n991, n992, n993, n994, n995, n996, n1061, n1062, n1063, 
        n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, 
        n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, 
        n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, 
        n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, 
        n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, 
        n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, 
        n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, 
        n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, 
        n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, 
        n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, 
        n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, 
        n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, 
        n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, 
        n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, 
        n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, 
        n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, 
        n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, 
        n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, 
        n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, 
        n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
        n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, 
        n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
        n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, 
        n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, 
        n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, 
        n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, 
        n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, 
        n1280, n1281, n1282, n1283, n1284, n1349, n1350, n1351, 
        n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, 
        n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, 
        n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
        n1376, n1377, n1378, n1379, n1380, n1416, n1421, n1423, 
        n1424, n1425, n1437, n1438, n1439, n1451, n1452, n1453, 
        n1465, n1466, n1467, n1479, n1480, n1481, n1493, n1494, 
        n1495, n1507, n1508, n1509, n1521, n1522, n1523, n1535, 
        n1536, n1537, n1549, n1550, n1551, n1563, n1564, n1565, 
        n1577, n1578, n1579, n1591, n1592, n1593, n1605, n1606, 
        n1607, n1619, n1620, n1621, n1633, n1634, n1635, n1647, 
        n1648, n1649, n1661, n1662, n1663, n1675, n1676, n1677, 
        n1689, n1690, n1691, n1703, n1704, n1705, n1717, n1718, 
        n1719, n1731, n1732, n1733, n1745, n1746, n1747, n1759, 
        n1760, n1761, n1773, n1774, n1775, n1787, n1788, n1789, 
        n1801, n1802, n1803, n1815, n1816, n1817, n1829, n1830, 
        n1831, n1843, n1844, n1845, n1857, n1858, n1859;
    
    assign func1_in[31] = func0_in[31];   // gpio_mux.v(15)
    assign func1_in[30] = func0_in[30];   // gpio_mux.v(15)
    assign func1_in[29] = func0_in[29];   // gpio_mux.v(15)
    assign func1_in[28] = func0_in[28];   // gpio_mux.v(15)
    assign func1_in[27] = func0_in[27];   // gpio_mux.v(15)
    assign func1_in[26] = func0_in[26];   // gpio_mux.v(15)
    assign func1_in[25] = func0_in[25];   // gpio_mux.v(15)
    assign func1_in[24] = func0_in[24];   // gpio_mux.v(15)
    assign func1_in[23] = func0_in[23];   // gpio_mux.v(15)
    assign func1_in[22] = func0_in[22];   // gpio_mux.v(15)
    assign func1_in[21] = func0_in[21];   // gpio_mux.v(15)
    assign func1_in[20] = func0_in[20];   // gpio_mux.v(15)
    assign func1_in[19] = func0_in[19];   // gpio_mux.v(15)
    assign func1_in[18] = func0_in[18];   // gpio_mux.v(15)
    assign func1_in[17] = func0_in[17];   // gpio_mux.v(15)
    assign func1_in[16] = func0_in[16];   // gpio_mux.v(15)
    assign func1_in[15] = func0_in[15];   // gpio_mux.v(15)
    assign func1_in[14] = func0_in[14];   // gpio_mux.v(15)
    assign func1_in[13] = func0_in[13];   // gpio_mux.v(15)
    assign func1_in[12] = func0_in[12];   // gpio_mux.v(15)
    assign func1_in[11] = func0_in[11];   // gpio_mux.v(15)
    assign func1_in[10] = func0_in[10];   // gpio_mux.v(15)
    assign func1_in[9] = func0_in[9];   // gpio_mux.v(15)
    assign func1_in[8] = func0_in[8];   // gpio_mux.v(15)
    assign func1_in[7] = func0_in[7];   // gpio_mux.v(15)
    assign func1_in[6] = func0_in[6];   // gpio_mux.v(15)
    assign func1_in[5] = func0_in[5];   // gpio_mux.v(15)
    assign func1_in[4] = func0_in[4];   // gpio_mux.v(15)
    assign func1_in[3] = func0_in[3];   // gpio_mux.v(15)
    assign func1_in[2] = func0_in[2];   // gpio_mux.v(15)
    assign func1_in[1] = func0_in[1];   // gpio_mux.v(15)
    assign func1_in[0] = func0_in[0];   // gpio_mux.v(15)
    assign func2_in[31] = func0_in[31];   // gpio_mux.v(16)
    assign func2_in[30] = func0_in[30];   // gpio_mux.v(16)
    assign func2_in[29] = func0_in[29];   // gpio_mux.v(16)
    assign func2_in[28] = func0_in[28];   // gpio_mux.v(16)
    assign func2_in[27] = func0_in[27];   // gpio_mux.v(16)
    assign func2_in[26] = func0_in[26];   // gpio_mux.v(16)
    assign func2_in[25] = func0_in[25];   // gpio_mux.v(16)
    assign func2_in[24] = func0_in[24];   // gpio_mux.v(16)
    assign func2_in[23] = func0_in[23];   // gpio_mux.v(16)
    assign func2_in[22] = func0_in[22];   // gpio_mux.v(16)
    assign func2_in[21] = func0_in[21];   // gpio_mux.v(16)
    assign func2_in[20] = func0_in[20];   // gpio_mux.v(16)
    assign func2_in[19] = func0_in[19];   // gpio_mux.v(16)
    assign func2_in[18] = func0_in[18];   // gpio_mux.v(16)
    assign func2_in[17] = func0_in[17];   // gpio_mux.v(16)
    assign func2_in[16] = func0_in[16];   // gpio_mux.v(16)
    assign func2_in[15] = func0_in[15];   // gpio_mux.v(16)
    assign func2_in[14] = func0_in[14];   // gpio_mux.v(16)
    assign func2_in[13] = func0_in[13];   // gpio_mux.v(16)
    assign func2_in[12] = func0_in[12];   // gpio_mux.v(16)
    assign func2_in[11] = func0_in[11];   // gpio_mux.v(16)
    assign func2_in[10] = func0_in[10];   // gpio_mux.v(16)
    assign func2_in[9] = func0_in[9];   // gpio_mux.v(16)
    assign func2_in[8] = func0_in[8];   // gpio_mux.v(16)
    assign func2_in[7] = func0_in[7];   // gpio_mux.v(16)
    assign func2_in[6] = func0_in[6];   // gpio_mux.v(16)
    assign func2_in[5] = func0_in[5];   // gpio_mux.v(16)
    assign func2_in[4] = func0_in[4];   // gpio_mux.v(16)
    assign func2_in[3] = func0_in[3];   // gpio_mux.v(16)
    assign func2_in[2] = func0_in[2];   // gpio_mux.v(16)
    assign func2_in[1] = func0_in[1];   // gpio_mux.v(16)
    assign func2_in[0] = func0_in[0];   // gpio_mux.v(16)
    assign func3_in[31] = func0_in[31];   // gpio_mux.v(17)
    assign func3_in[30] = func0_in[30];   // gpio_mux.v(17)
    assign func3_in[29] = func0_in[29];   // gpio_mux.v(17)
    assign func3_in[28] = func0_in[28];   // gpio_mux.v(17)
    assign func3_in[27] = func0_in[27];   // gpio_mux.v(17)
    assign func3_in[26] = func0_in[26];   // gpio_mux.v(17)
    assign func3_in[25] = func0_in[25];   // gpio_mux.v(17)
    assign func3_in[24] = func0_in[24];   // gpio_mux.v(17)
    assign func3_in[23] = func0_in[23];   // gpio_mux.v(17)
    assign func3_in[22] = func0_in[22];   // gpio_mux.v(17)
    assign func3_in[21] = func0_in[21];   // gpio_mux.v(17)
    assign func3_in[20] = func0_in[20];   // gpio_mux.v(17)
    assign func3_in[19] = func0_in[19];   // gpio_mux.v(17)
    assign func3_in[18] = func0_in[18];   // gpio_mux.v(17)
    assign func3_in[17] = func0_in[17];   // gpio_mux.v(17)
    assign func3_in[16] = func0_in[16];   // gpio_mux.v(17)
    assign func3_in[15] = func0_in[15];   // gpio_mux.v(17)
    assign func3_in[14] = func0_in[14];   // gpio_mux.v(17)
    assign func3_in[13] = func0_in[13];   // gpio_mux.v(17)
    assign func3_in[12] = func0_in[12];   // gpio_mux.v(17)
    assign func3_in[11] = func0_in[11];   // gpio_mux.v(17)
    assign func3_in[10] = func0_in[10];   // gpio_mux.v(17)
    assign func3_in[9] = func0_in[9];   // gpio_mux.v(17)
    assign func3_in[8] = func0_in[8];   // gpio_mux.v(17)
    assign func3_in[7] = func0_in[7];   // gpio_mux.v(17)
    assign func3_in[6] = func0_in[6];   // gpio_mux.v(17)
    assign func3_in[5] = func0_in[5];   // gpio_mux.v(17)
    assign func3_in[4] = func0_in[4];   // gpio_mux.v(17)
    assign func3_in[3] = func0_in[3];   // gpio_mux.v(17)
    assign func3_in[2] = func0_in[2];   // gpio_mux.v(17)
    assign func3_in[1] = func0_in[1];   // gpio_mux.v(17)
    assign func3_in[0] = func0_in[0];   // gpio_mux.v(17)
    nor (n4, \pin_mux[0].pin_control [1], \pin_mux[0].pin_control [0]) ;   // gpio_mux.v(48)
    not (n5, \pin_mux[0].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n6, \pin_mux[0].pin_control [1], n5) ;   // gpio_mux.v(48)
    not (n7, \pin_mux[0].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n8, n7, \pin_mux[0].pin_control [0]) ;   // gpio_mux.v(48)
    assign n9 = n8 ? func2_out[0] : func3_out[0];   // gpio_mux.v(48)
    assign n10 = n6 ? func1_out[0] : n9;   // gpio_mux.v(48)
    assign \pin_mux[0].pin_out  = n4 ? func0_out[0] : n10;   // gpio_mux.v(48)
    assign n17 = n8 ? func2_dir[0] : func3_dir[0];   // gpio_mux.v(49)
    assign n18 = n6 ? func1_dir[0] : n17;   // gpio_mux.v(49)
    assign \pin_mux[0].pin_dir  = n4 ? func0_dir[0] : n18;   // gpio_mux.v(49)
    assign pins[0] = \pin_mux[0].pin_dir  ? \pin_mux[0].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[0] = \pin_mux[0].pin_dir  ? \pin_mux[0].pin_out  : pins[0];   // gpio_mux.v(51)
    nor (n33, \pin_mux[1].pin_control [1], \pin_mux[1].pin_control [0]) ;   // gpio_mux.v(48)
    not (n34, \pin_mux[1].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n35, \pin_mux[1].pin_control [1], n34) ;   // gpio_mux.v(48)
    not (n36, \pin_mux[1].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n37, n36, \pin_mux[1].pin_control [0]) ;   // gpio_mux.v(48)
    assign n38 = n37 ? func2_out[1] : func3_out[1];   // gpio_mux.v(48)
    assign n39 = n35 ? func1_out[1] : n38;   // gpio_mux.v(48)
    assign \pin_mux[1].pin_out  = n33 ? func0_out[1] : n39;   // gpio_mux.v(48)
    assign n46 = n37 ? func2_dir[1] : func3_dir[1];   // gpio_mux.v(49)
    assign n47 = n35 ? func1_dir[1] : n46;   // gpio_mux.v(49)
    assign \pin_mux[1].pin_dir  = n33 ? func0_dir[1] : n47;   // gpio_mux.v(49)
    assign pins[1] = \pin_mux[1].pin_dir  ? \pin_mux[1].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[1] = \pin_mux[1].pin_dir  ? \pin_mux[1].pin_out  : pins[1];   // gpio_mux.v(51)
    nor (n62, \pin_mux[2].pin_control [1], \pin_mux[2].pin_control [0]) ;   // gpio_mux.v(48)
    not (n63, \pin_mux[2].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n64, \pin_mux[2].pin_control [1], n63) ;   // gpio_mux.v(48)
    not (n65, \pin_mux[2].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n66, n65, \pin_mux[2].pin_control [0]) ;   // gpio_mux.v(48)
    assign n67 = n66 ? func2_out[2] : func3_out[2];   // gpio_mux.v(48)
    assign n68 = n64 ? func1_out[2] : n67;   // gpio_mux.v(48)
    assign \pin_mux[2].pin_out  = n62 ? func0_out[2] : n68;   // gpio_mux.v(48)
    assign n75 = n66 ? func2_dir[2] : func3_dir[2];   // gpio_mux.v(49)
    assign n76 = n64 ? func1_dir[2] : n75;   // gpio_mux.v(49)
    assign \pin_mux[2].pin_dir  = n62 ? func0_dir[2] : n76;   // gpio_mux.v(49)
    assign pins[2] = \pin_mux[2].pin_dir  ? \pin_mux[2].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[2] = \pin_mux[2].pin_dir  ? \pin_mux[2].pin_out  : pins[2];   // gpio_mux.v(51)
    nor (n91, \pin_mux[3].pin_control [1], \pin_mux[3].pin_control [0]) ;   // gpio_mux.v(48)
    not (n92, \pin_mux[3].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n93, \pin_mux[3].pin_control [1], n92) ;   // gpio_mux.v(48)
    not (n94, \pin_mux[3].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n95, n94, \pin_mux[3].pin_control [0]) ;   // gpio_mux.v(48)
    assign n96 = n95 ? func2_out[3] : func3_out[3];   // gpio_mux.v(48)
    assign n97 = n93 ? func1_out[3] : n96;   // gpio_mux.v(48)
    assign \pin_mux[3].pin_out  = n91 ? func0_out[3] : n97;   // gpio_mux.v(48)
    assign n104 = n95 ? func2_dir[3] : func3_dir[3];   // gpio_mux.v(49)
    assign n105 = n93 ? func1_dir[3] : n104;   // gpio_mux.v(49)
    assign \pin_mux[3].pin_dir  = n91 ? func0_dir[3] : n105;   // gpio_mux.v(49)
    assign pins[3] = \pin_mux[3].pin_dir  ? \pin_mux[3].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[3] = \pin_mux[3].pin_dir  ? \pin_mux[3].pin_out  : pins[3];   // gpio_mux.v(51)
    nor (n120, \pin_mux[4].pin_control [1], \pin_mux[4].pin_control [0]) ;   // gpio_mux.v(48)
    not (n121, \pin_mux[4].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n122, \pin_mux[4].pin_control [1], n121) ;   // gpio_mux.v(48)
    not (n123, \pin_mux[4].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n124, n123, \pin_mux[4].pin_control [0]) ;   // gpio_mux.v(48)
    assign n125 = n124 ? func2_out[4] : func3_out[4];   // gpio_mux.v(48)
    assign n126 = n122 ? func1_out[4] : n125;   // gpio_mux.v(48)
    assign \pin_mux[4].pin_out  = n120 ? func0_out[4] : n126;   // gpio_mux.v(48)
    assign n133 = n124 ? func2_dir[4] : func3_dir[4];   // gpio_mux.v(49)
    assign n134 = n122 ? func1_dir[4] : n133;   // gpio_mux.v(49)
    assign \pin_mux[4].pin_dir  = n120 ? func0_dir[4] : n134;   // gpio_mux.v(49)
    assign pins[4] = \pin_mux[4].pin_dir  ? \pin_mux[4].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[4] = \pin_mux[4].pin_dir  ? \pin_mux[4].pin_out  : pins[4];   // gpio_mux.v(51)
    nor (n149, \pin_mux[5].pin_control [1], \pin_mux[5].pin_control [0]) ;   // gpio_mux.v(48)
    not (n150, \pin_mux[5].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n151, \pin_mux[5].pin_control [1], n150) ;   // gpio_mux.v(48)
    not (n152, \pin_mux[5].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n153, n152, \pin_mux[5].pin_control [0]) ;   // gpio_mux.v(48)
    assign n154 = n153 ? func2_out[5] : func3_out[5];   // gpio_mux.v(48)
    assign n155 = n151 ? func1_out[5] : n154;   // gpio_mux.v(48)
    assign \pin_mux[5].pin_out  = n149 ? func0_out[5] : n155;   // gpio_mux.v(48)
    assign n162 = n153 ? func2_dir[5] : func3_dir[5];   // gpio_mux.v(49)
    assign n163 = n151 ? func1_dir[5] : n162;   // gpio_mux.v(49)
    assign \pin_mux[5].pin_dir  = n149 ? func0_dir[5] : n163;   // gpio_mux.v(49)
    assign pins[5] = \pin_mux[5].pin_dir  ? \pin_mux[5].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[5] = \pin_mux[5].pin_dir  ? \pin_mux[5].pin_out  : pins[5];   // gpio_mux.v(51)
    nor (n178, \pin_mux[6].pin_control [1], \pin_mux[6].pin_control [0]) ;   // gpio_mux.v(48)
    not (n179, \pin_mux[6].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n180, \pin_mux[6].pin_control [1], n179) ;   // gpio_mux.v(48)
    not (n181, \pin_mux[6].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n182, n181, \pin_mux[6].pin_control [0]) ;   // gpio_mux.v(48)
    assign n183 = n182 ? func2_out[6] : func3_out[6];   // gpio_mux.v(48)
    assign n184 = n180 ? func1_out[6] : n183;   // gpio_mux.v(48)
    assign \pin_mux[6].pin_out  = n178 ? func0_out[6] : n184;   // gpio_mux.v(48)
    assign n191 = n182 ? func2_dir[6] : func3_dir[6];   // gpio_mux.v(49)
    assign n192 = n180 ? func1_dir[6] : n191;   // gpio_mux.v(49)
    assign \pin_mux[6].pin_dir  = n178 ? func0_dir[6] : n192;   // gpio_mux.v(49)
    assign pins[6] = \pin_mux[6].pin_dir  ? \pin_mux[6].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[6] = \pin_mux[6].pin_dir  ? \pin_mux[6].pin_out  : pins[6];   // gpio_mux.v(51)
    nor (n207, \pin_mux[7].pin_control [1], \pin_mux[7].pin_control [0]) ;   // gpio_mux.v(48)
    not (n208, \pin_mux[7].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n209, \pin_mux[7].pin_control [1], n208) ;   // gpio_mux.v(48)
    not (n210, \pin_mux[7].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n211, n210, \pin_mux[7].pin_control [0]) ;   // gpio_mux.v(48)
    assign n212 = n211 ? func2_out[7] : func3_out[7];   // gpio_mux.v(48)
    assign n213 = n209 ? func1_out[7] : n212;   // gpio_mux.v(48)
    assign \pin_mux[7].pin_out  = n207 ? func0_out[7] : n213;   // gpio_mux.v(48)
    assign n220 = n211 ? func2_dir[7] : func3_dir[7];   // gpio_mux.v(49)
    assign n221 = n209 ? func1_dir[7] : n220;   // gpio_mux.v(49)
    assign \pin_mux[7].pin_dir  = n207 ? func0_dir[7] : n221;   // gpio_mux.v(49)
    assign pins[7] = \pin_mux[7].pin_dir  ? \pin_mux[7].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[7] = \pin_mux[7].pin_dir  ? \pin_mux[7].pin_out  : pins[7];   // gpio_mux.v(51)
    nor (n236, \pin_mux[8].pin_control [1], \pin_mux[8].pin_control [0]) ;   // gpio_mux.v(48)
    not (n237, \pin_mux[8].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n238, \pin_mux[8].pin_control [1], n237) ;   // gpio_mux.v(48)
    not (n239, \pin_mux[8].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n240, n239, \pin_mux[8].pin_control [0]) ;   // gpio_mux.v(48)
    assign n241 = n240 ? func2_out[8] : func3_out[8];   // gpio_mux.v(48)
    assign n242 = n238 ? func1_out[8] : n241;   // gpio_mux.v(48)
    assign \pin_mux[8].pin_out  = n236 ? func0_out[8] : n242;   // gpio_mux.v(48)
    assign n249 = n240 ? func2_dir[8] : func3_dir[8];   // gpio_mux.v(49)
    assign n250 = n238 ? func1_dir[8] : n249;   // gpio_mux.v(49)
    assign \pin_mux[8].pin_dir  = n236 ? func0_dir[8] : n250;   // gpio_mux.v(49)
    assign pins[8] = \pin_mux[8].pin_dir  ? \pin_mux[8].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[8] = \pin_mux[8].pin_dir  ? \pin_mux[8].pin_out  : pins[8];   // gpio_mux.v(51)
    nor (n265, \pin_mux[9].pin_control [1], \pin_mux[9].pin_control [0]) ;   // gpio_mux.v(48)
    not (n266, \pin_mux[9].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n267, \pin_mux[9].pin_control [1], n266) ;   // gpio_mux.v(48)
    not (n268, \pin_mux[9].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n269, n268, \pin_mux[9].pin_control [0]) ;   // gpio_mux.v(48)
    assign n270 = n269 ? func2_out[9] : func3_out[9];   // gpio_mux.v(48)
    assign n271 = n267 ? func1_out[9] : n270;   // gpio_mux.v(48)
    assign \pin_mux[9].pin_out  = n265 ? func0_out[9] : n271;   // gpio_mux.v(48)
    assign n278 = n269 ? func2_dir[9] : func3_dir[9];   // gpio_mux.v(49)
    assign n279 = n267 ? func1_dir[9] : n278;   // gpio_mux.v(49)
    assign \pin_mux[9].pin_dir  = n265 ? func0_dir[9] : n279;   // gpio_mux.v(49)
    assign pins[9] = \pin_mux[9].pin_dir  ? \pin_mux[9].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[9] = \pin_mux[9].pin_dir  ? \pin_mux[9].pin_out  : pins[9];   // gpio_mux.v(51)
    nor (n294, \pin_mux[10].pin_control [1], \pin_mux[10].pin_control [0]) ;   // gpio_mux.v(48)
    not (n295, \pin_mux[10].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n296, \pin_mux[10].pin_control [1], n295) ;   // gpio_mux.v(48)
    not (n297, \pin_mux[10].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n298, n297, \pin_mux[10].pin_control [0]) ;   // gpio_mux.v(48)
    assign n299 = n298 ? func2_out[10] : func3_out[10];   // gpio_mux.v(48)
    assign n300 = n296 ? func1_out[10] : n299;   // gpio_mux.v(48)
    assign \pin_mux[10].pin_out  = n294 ? func0_out[10] : n300;   // gpio_mux.v(48)
    assign n307 = n298 ? func2_dir[10] : func3_dir[10];   // gpio_mux.v(49)
    assign n308 = n296 ? func1_dir[10] : n307;   // gpio_mux.v(49)
    assign \pin_mux[10].pin_dir  = n294 ? func0_dir[10] : n308;   // gpio_mux.v(49)
    assign pins[10] = \pin_mux[10].pin_dir  ? \pin_mux[10].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[10] = \pin_mux[10].pin_dir  ? \pin_mux[10].pin_out  : pins[10];   // gpio_mux.v(51)
    nor (n323, \pin_mux[11].pin_control [1], \pin_mux[11].pin_control [0]) ;   // gpio_mux.v(48)
    not (n324, \pin_mux[11].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n325, \pin_mux[11].pin_control [1], n324) ;   // gpio_mux.v(48)
    not (n326, \pin_mux[11].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n327, n326, \pin_mux[11].pin_control [0]) ;   // gpio_mux.v(48)
    assign n328 = n327 ? func2_out[11] : func3_out[11];   // gpio_mux.v(48)
    assign n329 = n325 ? func1_out[11] : n328;   // gpio_mux.v(48)
    assign \pin_mux[11].pin_out  = n323 ? func0_out[11] : n329;   // gpio_mux.v(48)
    assign n336 = n327 ? func2_dir[11] : func3_dir[11];   // gpio_mux.v(49)
    assign n337 = n325 ? func1_dir[11] : n336;   // gpio_mux.v(49)
    assign \pin_mux[11].pin_dir  = n323 ? func0_dir[11] : n337;   // gpio_mux.v(49)
    assign pins[11] = \pin_mux[11].pin_dir  ? \pin_mux[11].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[11] = \pin_mux[11].pin_dir  ? \pin_mux[11].pin_out  : pins[11];   // gpio_mux.v(51)
    nor (n352, \pin_mux[12].pin_control [1], \pin_mux[12].pin_control [0]) ;   // gpio_mux.v(48)
    not (n353, \pin_mux[12].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n354, \pin_mux[12].pin_control [1], n353) ;   // gpio_mux.v(48)
    not (n355, \pin_mux[12].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n356, n355, \pin_mux[12].pin_control [0]) ;   // gpio_mux.v(48)
    assign n357 = n356 ? func2_out[12] : func3_out[12];   // gpio_mux.v(48)
    assign n358 = n354 ? func1_out[12] : n357;   // gpio_mux.v(48)
    assign \pin_mux[12].pin_out  = n352 ? func0_out[12] : n358;   // gpio_mux.v(48)
    assign n365 = n356 ? func2_dir[12] : func3_dir[12];   // gpio_mux.v(49)
    assign n366 = n354 ? func1_dir[12] : n365;   // gpio_mux.v(49)
    assign \pin_mux[12].pin_dir  = n352 ? func0_dir[12] : n366;   // gpio_mux.v(49)
    assign pins[12] = \pin_mux[12].pin_dir  ? \pin_mux[12].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[12] = \pin_mux[12].pin_dir  ? \pin_mux[12].pin_out  : pins[12];   // gpio_mux.v(51)
    nor (n381, \pin_mux[13].pin_control [1], \pin_mux[13].pin_control [0]) ;   // gpio_mux.v(48)
    not (n382, \pin_mux[13].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n383, \pin_mux[13].pin_control [1], n382) ;   // gpio_mux.v(48)
    not (n384, \pin_mux[13].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n385, n384, \pin_mux[13].pin_control [0]) ;   // gpio_mux.v(48)
    assign n386 = n385 ? func2_out[13] : func3_out[13];   // gpio_mux.v(48)
    assign n387 = n383 ? func1_out[13] : n386;   // gpio_mux.v(48)
    assign \pin_mux[13].pin_out  = n381 ? func0_out[13] : n387;   // gpio_mux.v(48)
    assign n394 = n385 ? func2_dir[13] : func3_dir[13];   // gpio_mux.v(49)
    assign n395 = n383 ? func1_dir[13] : n394;   // gpio_mux.v(49)
    assign \pin_mux[13].pin_dir  = n381 ? func0_dir[13] : n395;   // gpio_mux.v(49)
    assign pins[13] = \pin_mux[13].pin_dir  ? \pin_mux[13].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[13] = \pin_mux[13].pin_dir  ? \pin_mux[13].pin_out  : pins[13];   // gpio_mux.v(51)
    nor (n410, \pin_mux[14].pin_control [1], \pin_mux[14].pin_control [0]) ;   // gpio_mux.v(48)
    not (n411, \pin_mux[14].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n412, \pin_mux[14].pin_control [1], n411) ;   // gpio_mux.v(48)
    not (n413, \pin_mux[14].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n414, n413, \pin_mux[14].pin_control [0]) ;   // gpio_mux.v(48)
    assign n415 = n414 ? func2_out[14] : func3_out[14];   // gpio_mux.v(48)
    assign n416 = n412 ? func1_out[14] : n415;   // gpio_mux.v(48)
    assign \pin_mux[14].pin_out  = n410 ? func0_out[14] : n416;   // gpio_mux.v(48)
    assign n423 = n414 ? func2_dir[14] : func3_dir[14];   // gpio_mux.v(49)
    assign n424 = n412 ? func1_dir[14] : n423;   // gpio_mux.v(49)
    assign \pin_mux[14].pin_dir  = n410 ? func0_dir[14] : n424;   // gpio_mux.v(49)
    assign pins[14] = \pin_mux[14].pin_dir  ? \pin_mux[14].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[14] = \pin_mux[14].pin_dir  ? \pin_mux[14].pin_out  : pins[14];   // gpio_mux.v(51)
    nor (n439, \pin_mux[15].pin_control [1], \pin_mux[15].pin_control [0]) ;   // gpio_mux.v(48)
    not (n440, \pin_mux[15].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n441, \pin_mux[15].pin_control [1], n440) ;   // gpio_mux.v(48)
    not (n442, \pin_mux[15].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n443, n442, \pin_mux[15].pin_control [0]) ;   // gpio_mux.v(48)
    assign n444 = n443 ? func2_out[15] : func3_out[15];   // gpio_mux.v(48)
    assign n445 = n441 ? func1_out[15] : n444;   // gpio_mux.v(48)
    assign \pin_mux[15].pin_out  = n439 ? func0_out[15] : n445;   // gpio_mux.v(48)
    assign n452 = n443 ? func2_dir[15] : func3_dir[15];   // gpio_mux.v(49)
    assign n453 = n441 ? func1_dir[15] : n452;   // gpio_mux.v(49)
    assign \pin_mux[15].pin_dir  = n439 ? func0_dir[15] : n453;   // gpio_mux.v(49)
    assign pins[15] = \pin_mux[15].pin_dir  ? \pin_mux[15].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[15] = \pin_mux[15].pin_dir  ? \pin_mux[15].pin_out  : pins[15];   // gpio_mux.v(51)
    nor (n468, \pin_mux[16].pin_control [1], \pin_mux[16].pin_control [0]) ;   // gpio_mux.v(48)
    not (n469, \pin_mux[16].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n470, \pin_mux[16].pin_control [1], n469) ;   // gpio_mux.v(48)
    not (n471, \pin_mux[16].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n472, n471, \pin_mux[16].pin_control [0]) ;   // gpio_mux.v(48)
    assign n473 = n472 ? func2_out[16] : func3_out[16];   // gpio_mux.v(48)
    assign n474 = n470 ? func1_out[16] : n473;   // gpio_mux.v(48)
    assign \pin_mux[16].pin_out  = n468 ? func0_out[16] : n474;   // gpio_mux.v(48)
    assign n481 = n472 ? func2_dir[16] : func3_dir[16];   // gpio_mux.v(49)
    assign n482 = n470 ? func1_dir[16] : n481;   // gpio_mux.v(49)
    assign \pin_mux[16].pin_dir  = n468 ? func0_dir[16] : n482;   // gpio_mux.v(49)
    assign pins[16] = \pin_mux[16].pin_dir  ? \pin_mux[16].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[16] = \pin_mux[16].pin_dir  ? \pin_mux[16].pin_out  : pins[16];   // gpio_mux.v(51)
    nor (n497, \pin_mux[17].pin_control [1], \pin_mux[17].pin_control [0]) ;   // gpio_mux.v(48)
    not (n498, \pin_mux[17].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n499, \pin_mux[17].pin_control [1], n498) ;   // gpio_mux.v(48)
    not (n500, \pin_mux[17].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n501, n500, \pin_mux[17].pin_control [0]) ;   // gpio_mux.v(48)
    assign n502 = n501 ? func2_out[17] : func3_out[17];   // gpio_mux.v(48)
    assign n503 = n499 ? func1_out[17] : n502;   // gpio_mux.v(48)
    assign \pin_mux[17].pin_out  = n497 ? func0_out[17] : n503;   // gpio_mux.v(48)
    assign n510 = n501 ? func2_dir[17] : func3_dir[17];   // gpio_mux.v(49)
    assign n511 = n499 ? func1_dir[17] : n510;   // gpio_mux.v(49)
    assign \pin_mux[17].pin_dir  = n497 ? func0_dir[17] : n511;   // gpio_mux.v(49)
    assign pins[17] = \pin_mux[17].pin_dir  ? \pin_mux[17].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[17] = \pin_mux[17].pin_dir  ? \pin_mux[17].pin_out  : pins[17];   // gpio_mux.v(51)
    nor (n526, \pin_mux[18].pin_control [1], \pin_mux[18].pin_control [0]) ;   // gpio_mux.v(48)
    not (n527, \pin_mux[18].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n528, \pin_mux[18].pin_control [1], n527) ;   // gpio_mux.v(48)
    not (n529, \pin_mux[18].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n530, n529, \pin_mux[18].pin_control [0]) ;   // gpio_mux.v(48)
    assign n531 = n530 ? func2_out[18] : func3_out[18];   // gpio_mux.v(48)
    assign n532 = n528 ? func1_out[18] : n531;   // gpio_mux.v(48)
    assign \pin_mux[18].pin_out  = n526 ? func0_out[18] : n532;   // gpio_mux.v(48)
    assign n539 = n530 ? func2_dir[18] : func3_dir[18];   // gpio_mux.v(49)
    assign n540 = n528 ? func1_dir[18] : n539;   // gpio_mux.v(49)
    assign \pin_mux[18].pin_dir  = n526 ? func0_dir[18] : n540;   // gpio_mux.v(49)
    assign pins[18] = \pin_mux[18].pin_dir  ? \pin_mux[18].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[18] = \pin_mux[18].pin_dir  ? \pin_mux[18].pin_out  : pins[18];   // gpio_mux.v(51)
    nor (n555, \pin_mux[19].pin_control [1], \pin_mux[19].pin_control [0]) ;   // gpio_mux.v(48)
    not (n556, \pin_mux[19].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n557, \pin_mux[19].pin_control [1], n556) ;   // gpio_mux.v(48)
    not (n558, \pin_mux[19].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n559, n558, \pin_mux[19].pin_control [0]) ;   // gpio_mux.v(48)
    assign n560 = n559 ? func2_out[19] : func3_out[19];   // gpio_mux.v(48)
    assign n561 = n557 ? func1_out[19] : n560;   // gpio_mux.v(48)
    assign \pin_mux[19].pin_out  = n555 ? func0_out[19] : n561;   // gpio_mux.v(48)
    assign n568 = n559 ? func2_dir[19] : func3_dir[19];   // gpio_mux.v(49)
    assign n569 = n557 ? func1_dir[19] : n568;   // gpio_mux.v(49)
    assign \pin_mux[19].pin_dir  = n555 ? func0_dir[19] : n569;   // gpio_mux.v(49)
    assign pins[19] = \pin_mux[19].pin_dir  ? \pin_mux[19].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[19] = \pin_mux[19].pin_dir  ? \pin_mux[19].pin_out  : pins[19];   // gpio_mux.v(51)
    nor (n584, \pin_mux[20].pin_control [1], \pin_mux[20].pin_control [0]) ;   // gpio_mux.v(48)
    not (n585, \pin_mux[20].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n586, \pin_mux[20].pin_control [1], n585) ;   // gpio_mux.v(48)
    not (n587, \pin_mux[20].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n588, n587, \pin_mux[20].pin_control [0]) ;   // gpio_mux.v(48)
    assign n589 = n588 ? func2_out[20] : func3_out[20];   // gpio_mux.v(48)
    assign n590 = n586 ? func1_out[20] : n589;   // gpio_mux.v(48)
    assign \pin_mux[20].pin_out  = n584 ? func0_out[20] : n590;   // gpio_mux.v(48)
    assign n597 = n588 ? func2_dir[20] : func3_dir[20];   // gpio_mux.v(49)
    assign n598 = n586 ? func1_dir[20] : n597;   // gpio_mux.v(49)
    assign \pin_mux[20].pin_dir  = n584 ? func0_dir[20] : n598;   // gpio_mux.v(49)
    assign pins[20] = \pin_mux[20].pin_dir  ? \pin_mux[20].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[20] = \pin_mux[20].pin_dir  ? \pin_mux[20].pin_out  : pins[20];   // gpio_mux.v(51)
    nor (n613, \pin_mux[21].pin_control [1], \pin_mux[21].pin_control [0]) ;   // gpio_mux.v(48)
    not (n614, \pin_mux[21].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n615, \pin_mux[21].pin_control [1], n614) ;   // gpio_mux.v(48)
    not (n616, \pin_mux[21].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n617, n616, \pin_mux[21].pin_control [0]) ;   // gpio_mux.v(48)
    assign n618 = n617 ? func2_out[21] : func3_out[21];   // gpio_mux.v(48)
    assign n619 = n615 ? func1_out[21] : n618;   // gpio_mux.v(48)
    assign \pin_mux[21].pin_out  = n613 ? func0_out[21] : n619;   // gpio_mux.v(48)
    assign n626 = n617 ? func2_dir[21] : func3_dir[21];   // gpio_mux.v(49)
    assign n627 = n615 ? func1_dir[21] : n626;   // gpio_mux.v(49)
    assign \pin_mux[21].pin_dir  = n613 ? func0_dir[21] : n627;   // gpio_mux.v(49)
    assign pins[21] = \pin_mux[21].pin_dir  ? \pin_mux[21].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[21] = \pin_mux[21].pin_dir  ? \pin_mux[21].pin_out  : pins[21];   // gpio_mux.v(51)
    nor (n642, \pin_mux[22].pin_control [1], \pin_mux[22].pin_control [0]) ;   // gpio_mux.v(48)
    not (n643, \pin_mux[22].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n644, \pin_mux[22].pin_control [1], n643) ;   // gpio_mux.v(48)
    not (n645, \pin_mux[22].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n646, n645, \pin_mux[22].pin_control [0]) ;   // gpio_mux.v(48)
    assign n647 = n646 ? func2_out[22] : func3_out[22];   // gpio_mux.v(48)
    assign n648 = n644 ? func1_out[22] : n647;   // gpio_mux.v(48)
    assign \pin_mux[22].pin_out  = n642 ? func0_out[22] : n648;   // gpio_mux.v(48)
    assign n655 = n646 ? func2_dir[22] : func3_dir[22];   // gpio_mux.v(49)
    assign n656 = n644 ? func1_dir[22] : n655;   // gpio_mux.v(49)
    assign \pin_mux[22].pin_dir  = n642 ? func0_dir[22] : n656;   // gpio_mux.v(49)
    assign pins[22] = \pin_mux[22].pin_dir  ? \pin_mux[22].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[22] = \pin_mux[22].pin_dir  ? \pin_mux[22].pin_out  : pins[22];   // gpio_mux.v(51)
    nor (n671, \pin_mux[23].pin_control [1], \pin_mux[23].pin_control [0]) ;   // gpio_mux.v(48)
    not (n672, \pin_mux[23].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n673, \pin_mux[23].pin_control [1], n672) ;   // gpio_mux.v(48)
    not (n674, \pin_mux[23].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n675, n674, \pin_mux[23].pin_control [0]) ;   // gpio_mux.v(48)
    assign n676 = n675 ? func2_out[23] : func3_out[23];   // gpio_mux.v(48)
    assign n677 = n673 ? func1_out[23] : n676;   // gpio_mux.v(48)
    assign \pin_mux[23].pin_out  = n671 ? func0_out[23] : n677;   // gpio_mux.v(48)
    assign n684 = n675 ? func2_dir[23] : func3_dir[23];   // gpio_mux.v(49)
    assign n685 = n673 ? func1_dir[23] : n684;   // gpio_mux.v(49)
    assign \pin_mux[23].pin_dir  = n671 ? func0_dir[23] : n685;   // gpio_mux.v(49)
    assign pins[23] = \pin_mux[23].pin_dir  ? \pin_mux[23].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[23] = \pin_mux[23].pin_dir  ? \pin_mux[23].pin_out  : pins[23];   // gpio_mux.v(51)
    nor (n700, \pin_mux[24].pin_control [1], \pin_mux[24].pin_control [0]) ;   // gpio_mux.v(48)
    not (n701, \pin_mux[24].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n702, \pin_mux[24].pin_control [1], n701) ;   // gpio_mux.v(48)
    not (n703, \pin_mux[24].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n704, n703, \pin_mux[24].pin_control [0]) ;   // gpio_mux.v(48)
    assign n705 = n704 ? func2_out[24] : func3_out[24];   // gpio_mux.v(48)
    assign n706 = n702 ? func1_out[24] : n705;   // gpio_mux.v(48)
    assign \pin_mux[24].pin_out  = n700 ? func0_out[24] : n706;   // gpio_mux.v(48)
    assign n713 = n704 ? func2_dir[24] : func3_dir[24];   // gpio_mux.v(49)
    assign n714 = n702 ? func1_dir[24] : n713;   // gpio_mux.v(49)
    assign \pin_mux[24].pin_dir  = n700 ? func0_dir[24] : n714;   // gpio_mux.v(49)
    assign pins[24] = \pin_mux[24].pin_dir  ? \pin_mux[24].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[24] = \pin_mux[24].pin_dir  ? \pin_mux[24].pin_out  : pins[24];   // gpio_mux.v(51)
    nor (n729, \pin_mux[25].pin_control [1], \pin_mux[25].pin_control [0]) ;   // gpio_mux.v(48)
    not (n730, \pin_mux[25].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n731, \pin_mux[25].pin_control [1], n730) ;   // gpio_mux.v(48)
    not (n732, \pin_mux[25].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n733, n732, \pin_mux[25].pin_control [0]) ;   // gpio_mux.v(48)
    assign n734 = n733 ? func2_out[25] : func3_out[25];   // gpio_mux.v(48)
    assign n735 = n731 ? func1_out[25] : n734;   // gpio_mux.v(48)
    assign \pin_mux[25].pin_out  = n729 ? func0_out[25] : n735;   // gpio_mux.v(48)
    assign n742 = n733 ? func2_dir[25] : func3_dir[25];   // gpio_mux.v(49)
    assign n743 = n731 ? func1_dir[25] : n742;   // gpio_mux.v(49)
    assign \pin_mux[25].pin_dir  = n729 ? func0_dir[25] : n743;   // gpio_mux.v(49)
    assign pins[25] = \pin_mux[25].pin_dir  ? \pin_mux[25].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[25] = \pin_mux[25].pin_dir  ? \pin_mux[25].pin_out  : pins[25];   // gpio_mux.v(51)
    nor (n758, \pin_mux[26].pin_control [1], \pin_mux[26].pin_control [0]) ;   // gpio_mux.v(48)
    not (n759, \pin_mux[26].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n760, \pin_mux[26].pin_control [1], n759) ;   // gpio_mux.v(48)
    not (n761, \pin_mux[26].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n762, n761, \pin_mux[26].pin_control [0]) ;   // gpio_mux.v(48)
    assign n763 = n762 ? func2_out[26] : func3_out[26];   // gpio_mux.v(48)
    assign n764 = n760 ? func1_out[26] : n763;   // gpio_mux.v(48)
    assign \pin_mux[26].pin_out  = n758 ? func0_out[26] : n764;   // gpio_mux.v(48)
    assign n771 = n762 ? func2_dir[26] : func3_dir[26];   // gpio_mux.v(49)
    assign n772 = n760 ? func1_dir[26] : n771;   // gpio_mux.v(49)
    assign \pin_mux[26].pin_dir  = n758 ? func0_dir[26] : n772;   // gpio_mux.v(49)
    assign pins[26] = \pin_mux[26].pin_dir  ? \pin_mux[26].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[26] = \pin_mux[26].pin_dir  ? \pin_mux[26].pin_out  : pins[26];   // gpio_mux.v(51)
    nor (n787, \pin_mux[27].pin_control [1], \pin_mux[27].pin_control [0]) ;   // gpio_mux.v(48)
    not (n788, \pin_mux[27].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n789, \pin_mux[27].pin_control [1], n788) ;   // gpio_mux.v(48)
    not (n790, \pin_mux[27].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n791, n790, \pin_mux[27].pin_control [0]) ;   // gpio_mux.v(48)
    assign n792 = n791 ? func2_out[27] : func3_out[27];   // gpio_mux.v(48)
    assign n793 = n789 ? func1_out[27] : n792;   // gpio_mux.v(48)
    assign \pin_mux[27].pin_out  = n787 ? func0_out[27] : n793;   // gpio_mux.v(48)
    assign n800 = n791 ? func2_dir[27] : func3_dir[27];   // gpio_mux.v(49)
    assign n801 = n789 ? func1_dir[27] : n800;   // gpio_mux.v(49)
    assign \pin_mux[27].pin_dir  = n787 ? func0_dir[27] : n801;   // gpio_mux.v(49)
    assign pins[27] = \pin_mux[27].pin_dir  ? \pin_mux[27].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[27] = \pin_mux[27].pin_dir  ? \pin_mux[27].pin_out  : pins[27];   // gpio_mux.v(51)
    nor (n816, \pin_mux[28].pin_control [1], \pin_mux[28].pin_control [0]) ;   // gpio_mux.v(48)
    not (n817, \pin_mux[28].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n818, \pin_mux[28].pin_control [1], n817) ;   // gpio_mux.v(48)
    not (n819, \pin_mux[28].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n820, n819, \pin_mux[28].pin_control [0]) ;   // gpio_mux.v(48)
    assign n821 = n820 ? func2_out[28] : func3_out[28];   // gpio_mux.v(48)
    assign n822 = n818 ? func1_out[28] : n821;   // gpio_mux.v(48)
    assign \pin_mux[28].pin_out  = n816 ? func0_out[28] : n822;   // gpio_mux.v(48)
    assign n829 = n820 ? func2_dir[28] : func3_dir[28];   // gpio_mux.v(49)
    assign n830 = n818 ? func1_dir[28] : n829;   // gpio_mux.v(49)
    assign \pin_mux[28].pin_dir  = n816 ? func0_dir[28] : n830;   // gpio_mux.v(49)
    assign pins[28] = \pin_mux[28].pin_dir  ? \pin_mux[28].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[28] = \pin_mux[28].pin_dir  ? \pin_mux[28].pin_out  : pins[28];   // gpio_mux.v(51)
    nor (n845, \pin_mux[29].pin_control [1], \pin_mux[29].pin_control [0]) ;   // gpio_mux.v(48)
    not (n846, \pin_mux[29].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n847, \pin_mux[29].pin_control [1], n846) ;   // gpio_mux.v(48)
    not (n848, \pin_mux[29].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n849, n848, \pin_mux[29].pin_control [0]) ;   // gpio_mux.v(48)
    assign n850 = n849 ? func2_out[29] : func3_out[29];   // gpio_mux.v(48)
    assign n851 = n847 ? func1_out[29] : n850;   // gpio_mux.v(48)
    assign \pin_mux[29].pin_out  = n845 ? func0_out[29] : n851;   // gpio_mux.v(48)
    assign n858 = n849 ? func2_dir[29] : func3_dir[29];   // gpio_mux.v(49)
    assign n859 = n847 ? func1_dir[29] : n858;   // gpio_mux.v(49)
    assign \pin_mux[29].pin_dir  = n845 ? func0_dir[29] : n859;   // gpio_mux.v(49)
    assign pins[29] = \pin_mux[29].pin_dir  ? \pin_mux[29].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[29] = \pin_mux[29].pin_dir  ? \pin_mux[29].pin_out  : pins[29];   // gpio_mux.v(51)
    nor (n874, \pin_mux[30].pin_control [1], \pin_mux[30].pin_control [0]) ;   // gpio_mux.v(48)
    not (n875, \pin_mux[30].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n876, \pin_mux[30].pin_control [1], n875) ;   // gpio_mux.v(48)
    not (n877, \pin_mux[30].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n878, n877, \pin_mux[30].pin_control [0]) ;   // gpio_mux.v(48)
    assign n879 = n878 ? func2_out[30] : func3_out[30];   // gpio_mux.v(48)
    assign n880 = n876 ? func1_out[30] : n879;   // gpio_mux.v(48)
    assign \pin_mux[30].pin_out  = n874 ? func0_out[30] : n880;   // gpio_mux.v(48)
    assign n887 = n878 ? func2_dir[30] : func3_dir[30];   // gpio_mux.v(49)
    assign n888 = n876 ? func1_dir[30] : n887;   // gpio_mux.v(49)
    assign \pin_mux[30].pin_dir  = n874 ? func0_dir[30] : n888;   // gpio_mux.v(49)
    assign pins[30] = \pin_mux[30].pin_dir  ? \pin_mux[30].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[30] = \pin_mux[30].pin_dir  ? \pin_mux[30].pin_out  : pins[30];   // gpio_mux.v(51)
    nor (n903, \pin_mux[31].pin_control [1], \pin_mux[31].pin_control [0]) ;   // gpio_mux.v(48)
    not (n904, \pin_mux[31].pin_control [0]) ;   // gpio_mux.v(48)
    nor (n905, \pin_mux[31].pin_control [1], n904) ;   // gpio_mux.v(48)
    not (n906, \pin_mux[31].pin_control [1]) ;   // gpio_mux.v(48)
    nor (n907, n906, \pin_mux[31].pin_control [0]) ;   // gpio_mux.v(48)
    assign n908 = n907 ? func2_out[31] : func3_out[31];   // gpio_mux.v(48)
    assign n909 = n905 ? func1_out[31] : n908;   // gpio_mux.v(48)
    assign \pin_mux[31].pin_out  = n903 ? func0_out[31] : n909;   // gpio_mux.v(48)
    assign n916 = n907 ? func2_dir[31] : func3_dir[31];   // gpio_mux.v(49)
    assign n917 = n905 ? func1_dir[31] : n916;   // gpio_mux.v(49)
    assign \pin_mux[31].pin_dir  = n903 ? func0_dir[31] : n917;   // gpio_mux.v(49)
    assign pins[31] = \pin_mux[31].pin_dir  ? \pin_mux[31].pin_out  : 1'bz;   // gpio_mux.v(50)
    assign func0_in[31] = \pin_mux[31].pin_dir  ? \pin_mux[31].pin_out  : pins[31];   // gpio_mux.v(51)
    xor (n933, sys_r_addr[1], addr[1]) ;   // gpio_mux.v(65)
    xor (n934, sys_r_addr[2], addr[2]) ;   // gpio_mux.v(65)
    xor (n935, sys_r_addr[3], addr[3]) ;   // gpio_mux.v(65)
    xor (n936, sys_r_addr[4], addr[4]) ;   // gpio_mux.v(65)
    xor (n937, sys_r_addr[5], addr[5]) ;   // gpio_mux.v(65)
    xor (n938, sys_r_addr[6], addr[6]) ;   // gpio_mux.v(65)
    xor (n939, sys_r_addr[7], addr[7]) ;   // gpio_mux.v(65)
    xor (n940, sys_r_addr[8], addr[8]) ;   // gpio_mux.v(65)
    xor (n941, sys_r_addr[9], addr[9]) ;   // gpio_mux.v(65)
    xor (n942, sys_r_addr[10], addr[10]) ;   // gpio_mux.v(65)
    xor (n943, sys_r_addr[11], addr[11]) ;   // gpio_mux.v(65)
    xor (n944, sys_r_addr[12], addr[12]) ;   // gpio_mux.v(65)
    xor (n945, sys_r_addr[13], addr[13]) ;   // gpio_mux.v(65)
    xor (n946, sys_r_addr[14], addr[14]) ;   // gpio_mux.v(65)
    xor (n947, sys_r_addr[15], addr[15]) ;   // gpio_mux.v(65)
    xor (n948, sys_r_addr[16], addr[16]) ;   // gpio_mux.v(65)
    xor (n949, sys_r_addr[17], addr[17]) ;   // gpio_mux.v(65)
    xor (n950, sys_r_addr[18], addr[18]) ;   // gpio_mux.v(65)
    xor (n951, sys_r_addr[19], addr[19]) ;   // gpio_mux.v(65)
    xor (n952, sys_r_addr[20], addr[20]) ;   // gpio_mux.v(65)
    xor (n953, sys_r_addr[21], addr[21]) ;   // gpio_mux.v(65)
    xor (n954, sys_r_addr[22], addr[22]) ;   // gpio_mux.v(65)
    xor (n955, sys_r_addr[23], addr[23]) ;   // gpio_mux.v(65)
    xor (n956, sys_r_addr[24], addr[24]) ;   // gpio_mux.v(65)
    xor (n957, sys_r_addr[25], addr[25]) ;   // gpio_mux.v(65)
    xor (n958, sys_r_addr[26], addr[26]) ;   // gpio_mux.v(65)
    xor (n959, sys_r_addr[27], addr[27]) ;   // gpio_mux.v(65)
    xor (n960, sys_r_addr[28], addr[28]) ;   // gpio_mux.v(65)
    xor (n961, sys_r_addr[29], addr[29]) ;   // gpio_mux.v(65)
    xor (n962, sys_r_addr[30], addr[30]) ;   // gpio_mux.v(65)
    xor (n963, sys_r_addr[31], addr[31]) ;   // gpio_mux.v(65)
    nor (n964, n963, n962, n961, n960, n959, n958, n957, n956, 
        n955, n954, n953, n952, n951, n950, n949, n948, n947, 
        n946, n945, n944, n943, n942, n941, n940, n939, n938, 
        n937, n936, n935, n934, n933) ;   // gpio_mux.v(65)
    assign n965 = sys_r_addr[0] ? \pin_mux[31].pin_control [1] : \pin_mux[15].pin_control [1];   // gpio_mux.v(68)
    assign n966 = sys_r_addr[0] ? \pin_mux[31].pin_control [0] : \pin_mux[15].pin_control [0];   // gpio_mux.v(68)
    assign n967 = sys_r_addr[0] ? \pin_mux[30].pin_control [1] : \pin_mux[14].pin_control [1];   // gpio_mux.v(68)
    assign n968 = sys_r_addr[0] ? \pin_mux[30].pin_control [0] : \pin_mux[14].pin_control [0];   // gpio_mux.v(68)
    assign n969 = sys_r_addr[0] ? \pin_mux[29].pin_control [1] : \pin_mux[13].pin_control [1];   // gpio_mux.v(68)
    assign n970 = sys_r_addr[0] ? \pin_mux[29].pin_control [0] : \pin_mux[13].pin_control [0];   // gpio_mux.v(68)
    assign n971 = sys_r_addr[0] ? \pin_mux[28].pin_control [1] : \pin_mux[12].pin_control [1];   // gpio_mux.v(68)
    assign n972 = sys_r_addr[0] ? \pin_mux[28].pin_control [0] : \pin_mux[12].pin_control [0];   // gpio_mux.v(68)
    assign n973 = sys_r_addr[0] ? \pin_mux[27].pin_control [1] : \pin_mux[11].pin_control [1];   // gpio_mux.v(68)
    assign n974 = sys_r_addr[0] ? \pin_mux[27].pin_control [0] : \pin_mux[11].pin_control [0];   // gpio_mux.v(68)
    assign n975 = sys_r_addr[0] ? \pin_mux[26].pin_control [1] : \pin_mux[10].pin_control [1];   // gpio_mux.v(68)
    assign n976 = sys_r_addr[0] ? \pin_mux[26].pin_control [0] : \pin_mux[10].pin_control [0];   // gpio_mux.v(68)
    assign n977 = sys_r_addr[0] ? \pin_mux[25].pin_control [1] : \pin_mux[9].pin_control [1];   // gpio_mux.v(68)
    assign n978 = sys_r_addr[0] ? \pin_mux[25].pin_control [0] : \pin_mux[9].pin_control [0];   // gpio_mux.v(68)
    assign n979 = sys_r_addr[0] ? \pin_mux[24].pin_control [1] : \pin_mux[8].pin_control [1];   // gpio_mux.v(68)
    assign n980 = sys_r_addr[0] ? \pin_mux[24].pin_control [0] : \pin_mux[8].pin_control [0];   // gpio_mux.v(68)
    assign n981 = sys_r_addr[0] ? \pin_mux[23].pin_control [1] : \pin_mux[7].pin_control [1];   // gpio_mux.v(68)
    assign n982 = sys_r_addr[0] ? \pin_mux[23].pin_control [0] : \pin_mux[7].pin_control [0];   // gpio_mux.v(68)
    assign n983 = sys_r_addr[0] ? \pin_mux[22].pin_control [1] : \pin_mux[6].pin_control [1];   // gpio_mux.v(68)
    assign n984 = sys_r_addr[0] ? \pin_mux[22].pin_control [0] : \pin_mux[6].pin_control [0];   // gpio_mux.v(68)
    assign n985 = sys_r_addr[0] ? \pin_mux[21].pin_control [1] : \pin_mux[5].pin_control [1];   // gpio_mux.v(68)
    assign n986 = sys_r_addr[0] ? \pin_mux[21].pin_control [0] : \pin_mux[5].pin_control [0];   // gpio_mux.v(68)
    assign n987 = sys_r_addr[0] ? \pin_mux[20].pin_control [1] : \pin_mux[4].pin_control [1];   // gpio_mux.v(68)
    assign n988 = sys_r_addr[0] ? \pin_mux[20].pin_control [0] : \pin_mux[4].pin_control [0];   // gpio_mux.v(68)
    assign n989 = sys_r_addr[0] ? \pin_mux[19].pin_control [1] : \pin_mux[3].pin_control [1];   // gpio_mux.v(68)
    assign n990 = sys_r_addr[0] ? \pin_mux[19].pin_control [0] : \pin_mux[3].pin_control [0];   // gpio_mux.v(68)
    assign n991 = sys_r_addr[0] ? \pin_mux[18].pin_control [1] : \pin_mux[2].pin_control [1];   // gpio_mux.v(68)
    assign n992 = sys_r_addr[0] ? \pin_mux[18].pin_control [0] : \pin_mux[2].pin_control [0];   // gpio_mux.v(68)
    assign n993 = sys_r_addr[0] ? \pin_mux[17].pin_control [1] : \pin_mux[1].pin_control [1];   // gpio_mux.v(68)
    assign n994 = sys_r_addr[0] ? \pin_mux[17].pin_control [0] : \pin_mux[1].pin_control [0];   // gpio_mux.v(68)
    assign n995 = sys_r_addr[0] ? \pin_mux[16].pin_control [1] : \pin_mux[0].pin_control [1];   // gpio_mux.v(68)
    assign n996 = sys_r_addr[0] ? \pin_mux[16].pin_control [0] : \pin_mux[0].pin_control [0];   // gpio_mux.v(68)
    xor (n1061, sys_w_addr[1], addr[1]) ;   // gpio_mux.v(78)
    xor (n1062, sys_w_addr[2], addr[2]) ;   // gpio_mux.v(78)
    xor (n1063, sys_w_addr[3], addr[3]) ;   // gpio_mux.v(78)
    xor (n1064, sys_w_addr[4], addr[4]) ;   // gpio_mux.v(78)
    xor (n1065, sys_w_addr[5], addr[5]) ;   // gpio_mux.v(78)
    xor (n1066, sys_w_addr[6], addr[6]) ;   // gpio_mux.v(78)
    xor (n1067, sys_w_addr[7], addr[7]) ;   // gpio_mux.v(78)
    xor (n1068, sys_w_addr[8], addr[8]) ;   // gpio_mux.v(78)
    xor (n1069, sys_w_addr[9], addr[9]) ;   // gpio_mux.v(78)
    xor (n1070, sys_w_addr[10], addr[10]) ;   // gpio_mux.v(78)
    xor (n1071, sys_w_addr[11], addr[11]) ;   // gpio_mux.v(78)
    xor (n1072, sys_w_addr[12], addr[12]) ;   // gpio_mux.v(78)
    xor (n1073, sys_w_addr[13], addr[13]) ;   // gpio_mux.v(78)
    xor (n1074, sys_w_addr[14], addr[14]) ;   // gpio_mux.v(78)
    xor (n1075, sys_w_addr[15], addr[15]) ;   // gpio_mux.v(78)
    xor (n1076, sys_w_addr[16], addr[16]) ;   // gpio_mux.v(78)
    xor (n1077, sys_w_addr[17], addr[17]) ;   // gpio_mux.v(78)
    xor (n1078, sys_w_addr[18], addr[18]) ;   // gpio_mux.v(78)
    xor (n1079, sys_w_addr[19], addr[19]) ;   // gpio_mux.v(78)
    xor (n1080, sys_w_addr[20], addr[20]) ;   // gpio_mux.v(78)
    xor (n1081, sys_w_addr[21], addr[21]) ;   // gpio_mux.v(78)
    xor (n1082, sys_w_addr[22], addr[22]) ;   // gpio_mux.v(78)
    xor (n1083, sys_w_addr[23], addr[23]) ;   // gpio_mux.v(78)
    xor (n1084, sys_w_addr[24], addr[24]) ;   // gpio_mux.v(78)
    xor (n1085, sys_w_addr[25], addr[25]) ;   // gpio_mux.v(78)
    xor (n1086, sys_w_addr[26], addr[26]) ;   // gpio_mux.v(78)
    xor (n1087, sys_w_addr[27], addr[27]) ;   // gpio_mux.v(78)
    xor (n1088, sys_w_addr[28], addr[28]) ;   // gpio_mux.v(78)
    xor (n1089, sys_w_addr[29], addr[29]) ;   // gpio_mux.v(78)
    xor (n1090, sys_w_addr[30], addr[30]) ;   // gpio_mux.v(78)
    xor (n1091, sys_w_addr[31], addr[31]) ;   // gpio_mux.v(78)
    nor (n1092, n1091, n1090, n1089, n1088, n1087, n1086, n1085, 
        n1084, n1083, n1082, n1081, n1080, n1079, n1078, n1077, 
        n1076, n1075, n1074, n1073, n1072, n1071, n1070, n1069, 
        n1068, n1067, n1066, n1065, n1064, n1063, n1062, n1061) ;   // gpio_mux.v(78)
    assign n1093 = sys_w_addr[0] ? sys_w_line[31] : \pin_mux[31].pin_control [1];   // gpio_mux.v(81)
    assign n1094 = sys_w_addr[0] ? sys_w_line[30] : \pin_mux[31].pin_control [0];   // gpio_mux.v(81)
    assign n1095 = sys_w_addr[0] ? sys_w_line[29] : \pin_mux[30].pin_control [1];   // gpio_mux.v(81)
    assign n1096 = sys_w_addr[0] ? sys_w_line[28] : \pin_mux[30].pin_control [0];   // gpio_mux.v(81)
    assign n1097 = sys_w_addr[0] ? sys_w_line[27] : \pin_mux[29].pin_control [1];   // gpio_mux.v(81)
    assign n1098 = sys_w_addr[0] ? sys_w_line[26] : \pin_mux[29].pin_control [0];   // gpio_mux.v(81)
    assign n1099 = sys_w_addr[0] ? sys_w_line[25] : \pin_mux[28].pin_control [1];   // gpio_mux.v(81)
    assign n1100 = sys_w_addr[0] ? sys_w_line[24] : \pin_mux[28].pin_control [0];   // gpio_mux.v(81)
    assign n1101 = sys_w_addr[0] ? sys_w_line[23] : \pin_mux[27].pin_control [1];   // gpio_mux.v(81)
    assign n1102 = sys_w_addr[0] ? sys_w_line[22] : \pin_mux[27].pin_control [0];   // gpio_mux.v(81)
    assign n1103 = sys_w_addr[0] ? sys_w_line[21] : \pin_mux[26].pin_control [1];   // gpio_mux.v(81)
    assign n1104 = sys_w_addr[0] ? sys_w_line[20] : \pin_mux[26].pin_control [0];   // gpio_mux.v(81)
    assign n1105 = sys_w_addr[0] ? sys_w_line[19] : \pin_mux[25].pin_control [1];   // gpio_mux.v(81)
    assign n1106 = sys_w_addr[0] ? sys_w_line[18] : \pin_mux[25].pin_control [0];   // gpio_mux.v(81)
    assign n1107 = sys_w_addr[0] ? sys_w_line[17] : \pin_mux[24].pin_control [1];   // gpio_mux.v(81)
    assign n1108 = sys_w_addr[0] ? sys_w_line[16] : \pin_mux[24].pin_control [0];   // gpio_mux.v(81)
    assign n1109 = sys_w_addr[0] ? sys_w_line[15] : \pin_mux[23].pin_control [1];   // gpio_mux.v(81)
    assign n1110 = sys_w_addr[0] ? sys_w_line[14] : \pin_mux[23].pin_control [0];   // gpio_mux.v(81)
    assign n1111 = sys_w_addr[0] ? sys_w_line[13] : \pin_mux[22].pin_control [1];   // gpio_mux.v(81)
    assign n1112 = sys_w_addr[0] ? sys_w_line[12] : \pin_mux[22].pin_control [0];   // gpio_mux.v(81)
    assign n1113 = sys_w_addr[0] ? sys_w_line[11] : \pin_mux[21].pin_control [1];   // gpio_mux.v(81)
    assign n1114 = sys_w_addr[0] ? sys_w_line[10] : \pin_mux[21].pin_control [0];   // gpio_mux.v(81)
    assign n1115 = sys_w_addr[0] ? sys_w_line[9] : \pin_mux[20].pin_control [1];   // gpio_mux.v(81)
    assign n1116 = sys_w_addr[0] ? sys_w_line[8] : \pin_mux[20].pin_control [0];   // gpio_mux.v(81)
    assign n1117 = sys_w_addr[0] ? sys_w_line[7] : \pin_mux[19].pin_control [1];   // gpio_mux.v(81)
    assign n1118 = sys_w_addr[0] ? sys_w_line[6] : \pin_mux[19].pin_control [0];   // gpio_mux.v(81)
    assign n1119 = sys_w_addr[0] ? sys_w_line[5] : \pin_mux[18].pin_control [1];   // gpio_mux.v(81)
    assign n1120 = sys_w_addr[0] ? sys_w_line[4] : \pin_mux[18].pin_control [0];   // gpio_mux.v(81)
    assign n1121 = sys_w_addr[0] ? sys_w_line[3] : \pin_mux[17].pin_control [1];   // gpio_mux.v(81)
    assign n1122 = sys_w_addr[0] ? sys_w_line[2] : \pin_mux[17].pin_control [0];   // gpio_mux.v(81)
    assign n1123 = sys_w_addr[0] ? sys_w_line[1] : \pin_mux[16].pin_control [1];   // gpio_mux.v(81)
    assign n1124 = sys_w_addr[0] ? sys_w_line[0] : \pin_mux[16].pin_control [0];   // gpio_mux.v(81)
    assign n1125 = sys_w_addr[0] ? \pin_mux[15].pin_control [1] : sys_w_line[31];   // gpio_mux.v(81)
    assign n1126 = sys_w_addr[0] ? \pin_mux[15].pin_control [0] : sys_w_line[30];   // gpio_mux.v(81)
    assign n1127 = sys_w_addr[0] ? \pin_mux[14].pin_control [1] : sys_w_line[29];   // gpio_mux.v(81)
    assign n1128 = sys_w_addr[0] ? \pin_mux[14].pin_control [0] : sys_w_line[28];   // gpio_mux.v(81)
    assign n1129 = sys_w_addr[0] ? \pin_mux[13].pin_control [1] : sys_w_line[27];   // gpio_mux.v(81)
    assign n1130 = sys_w_addr[0] ? \pin_mux[13].pin_control [0] : sys_w_line[26];   // gpio_mux.v(81)
    assign n1131 = sys_w_addr[0] ? \pin_mux[12].pin_control [1] : sys_w_line[25];   // gpio_mux.v(81)
    assign n1132 = sys_w_addr[0] ? \pin_mux[12].pin_control [0] : sys_w_line[24];   // gpio_mux.v(81)
    assign n1133 = sys_w_addr[0] ? \pin_mux[11].pin_control [1] : sys_w_line[23];   // gpio_mux.v(81)
    assign n1134 = sys_w_addr[0] ? \pin_mux[11].pin_control [0] : sys_w_line[22];   // gpio_mux.v(81)
    assign n1135 = sys_w_addr[0] ? \pin_mux[10].pin_control [1] : sys_w_line[21];   // gpio_mux.v(81)
    assign n1136 = sys_w_addr[0] ? \pin_mux[10].pin_control [0] : sys_w_line[20];   // gpio_mux.v(81)
    assign n1137 = sys_w_addr[0] ? \pin_mux[9].pin_control [1] : sys_w_line[19];   // gpio_mux.v(81)
    assign n1138 = sys_w_addr[0] ? \pin_mux[9].pin_control [0] : sys_w_line[18];   // gpio_mux.v(81)
    assign n1139 = sys_w_addr[0] ? \pin_mux[8].pin_control [1] : sys_w_line[17];   // gpio_mux.v(81)
    assign n1140 = sys_w_addr[0] ? \pin_mux[8].pin_control [0] : sys_w_line[16];   // gpio_mux.v(81)
    assign n1141 = sys_w_addr[0] ? \pin_mux[7].pin_control [1] : sys_w_line[15];   // gpio_mux.v(81)
    assign n1142 = sys_w_addr[0] ? \pin_mux[7].pin_control [0] : sys_w_line[14];   // gpio_mux.v(81)
    assign n1143 = sys_w_addr[0] ? \pin_mux[6].pin_control [1] : sys_w_line[13];   // gpio_mux.v(81)
    assign n1144 = sys_w_addr[0] ? \pin_mux[6].pin_control [0] : sys_w_line[12];   // gpio_mux.v(81)
    assign n1145 = sys_w_addr[0] ? \pin_mux[5].pin_control [1] : sys_w_line[11];   // gpio_mux.v(81)
    assign n1146 = sys_w_addr[0] ? \pin_mux[5].pin_control [0] : sys_w_line[10];   // gpio_mux.v(81)
    assign n1147 = sys_w_addr[0] ? \pin_mux[4].pin_control [1] : sys_w_line[9];   // gpio_mux.v(81)
    assign n1148 = sys_w_addr[0] ? \pin_mux[4].pin_control [0] : sys_w_line[8];   // gpio_mux.v(81)
    assign n1149 = sys_w_addr[0] ? \pin_mux[3].pin_control [1] : sys_w_line[7];   // gpio_mux.v(81)
    assign n1150 = sys_w_addr[0] ? \pin_mux[3].pin_control [0] : sys_w_line[6];   // gpio_mux.v(81)
    assign n1151 = sys_w_addr[0] ? \pin_mux[2].pin_control [1] : sys_w_line[5];   // gpio_mux.v(81)
    assign n1152 = sys_w_addr[0] ? \pin_mux[2].pin_control [0] : sys_w_line[4];   // gpio_mux.v(81)
    assign n1153 = sys_w_addr[0] ? \pin_mux[1].pin_control [1] : sys_w_line[3];   // gpio_mux.v(81)
    assign n1154 = sys_w_addr[0] ? \pin_mux[1].pin_control [0] : sys_w_line[2];   // gpio_mux.v(81)
    assign n1155 = sys_w_addr[0] ? \pin_mux[0].pin_control [1] : sys_w_line[1];   // gpio_mux.v(81)
    assign n1156 = sys_w_addr[0] ? \pin_mux[0].pin_control [0] : sys_w_line[0];   // gpio_mux.v(81)
    assign n1157 = n1092 ? n1093 : \pin_mux[31].pin_control [1];   // gpio_mux.v(78)
    assign n1158 = n1092 ? n1094 : \pin_mux[31].pin_control [0];   // gpio_mux.v(78)
    assign n1159 = n1092 ? n1095 : \pin_mux[30].pin_control [1];   // gpio_mux.v(78)
    assign n1160 = n1092 ? n1096 : \pin_mux[30].pin_control [0];   // gpio_mux.v(78)
    assign n1161 = n1092 ? n1097 : \pin_mux[29].pin_control [1];   // gpio_mux.v(78)
    assign n1162 = n1092 ? n1098 : \pin_mux[29].pin_control [0];   // gpio_mux.v(78)
    assign n1163 = n1092 ? n1099 : \pin_mux[28].pin_control [1];   // gpio_mux.v(78)
    assign n1164 = n1092 ? n1100 : \pin_mux[28].pin_control [0];   // gpio_mux.v(78)
    assign n1165 = n1092 ? n1101 : \pin_mux[27].pin_control [1];   // gpio_mux.v(78)
    assign n1166 = n1092 ? n1102 : \pin_mux[27].pin_control [0];   // gpio_mux.v(78)
    assign n1167 = n1092 ? n1103 : \pin_mux[26].pin_control [1];   // gpio_mux.v(78)
    assign n1168 = n1092 ? n1104 : \pin_mux[26].pin_control [0];   // gpio_mux.v(78)
    assign n1169 = n1092 ? n1105 : \pin_mux[25].pin_control [1];   // gpio_mux.v(78)
    assign n1170 = n1092 ? n1106 : \pin_mux[25].pin_control [0];   // gpio_mux.v(78)
    assign n1171 = n1092 ? n1107 : \pin_mux[24].pin_control [1];   // gpio_mux.v(78)
    assign n1172 = n1092 ? n1108 : \pin_mux[24].pin_control [0];   // gpio_mux.v(78)
    assign n1173 = n1092 ? n1109 : \pin_mux[23].pin_control [1];   // gpio_mux.v(78)
    assign n1174 = n1092 ? n1110 : \pin_mux[23].pin_control [0];   // gpio_mux.v(78)
    assign n1175 = n1092 ? n1111 : \pin_mux[22].pin_control [1];   // gpio_mux.v(78)
    assign n1176 = n1092 ? n1112 : \pin_mux[22].pin_control [0];   // gpio_mux.v(78)
    assign n1177 = n1092 ? n1113 : \pin_mux[21].pin_control [1];   // gpio_mux.v(78)
    assign n1178 = n1092 ? n1114 : \pin_mux[21].pin_control [0];   // gpio_mux.v(78)
    assign n1179 = n1092 ? n1115 : \pin_mux[20].pin_control [1];   // gpio_mux.v(78)
    assign n1180 = n1092 ? n1116 : \pin_mux[20].pin_control [0];   // gpio_mux.v(78)
    assign n1181 = n1092 ? n1117 : \pin_mux[19].pin_control [1];   // gpio_mux.v(78)
    assign n1182 = n1092 ? n1118 : \pin_mux[19].pin_control [0];   // gpio_mux.v(78)
    assign n1183 = n1092 ? n1119 : \pin_mux[18].pin_control [1];   // gpio_mux.v(78)
    assign n1184 = n1092 ? n1120 : \pin_mux[18].pin_control [0];   // gpio_mux.v(78)
    assign n1185 = n1092 ? n1121 : \pin_mux[17].pin_control [1];   // gpio_mux.v(78)
    assign n1186 = n1092 ? n1122 : \pin_mux[17].pin_control [0];   // gpio_mux.v(78)
    assign n1187 = n1092 ? n1123 : \pin_mux[16].pin_control [1];   // gpio_mux.v(78)
    assign n1188 = n1092 ? n1124 : \pin_mux[16].pin_control [0];   // gpio_mux.v(78)
    assign n1189 = n1092 ? n1125 : \pin_mux[15].pin_control [1];   // gpio_mux.v(78)
    assign n1190 = n1092 ? n1126 : \pin_mux[15].pin_control [0];   // gpio_mux.v(78)
    assign n1191 = n1092 ? n1127 : \pin_mux[14].pin_control [1];   // gpio_mux.v(78)
    assign n1192 = n1092 ? n1128 : \pin_mux[14].pin_control [0];   // gpio_mux.v(78)
    assign n1193 = n1092 ? n1129 : \pin_mux[13].pin_control [1];   // gpio_mux.v(78)
    assign n1194 = n1092 ? n1130 : \pin_mux[13].pin_control [0];   // gpio_mux.v(78)
    assign n1195 = n1092 ? n1131 : \pin_mux[12].pin_control [1];   // gpio_mux.v(78)
    assign n1196 = n1092 ? n1132 : \pin_mux[12].pin_control [0];   // gpio_mux.v(78)
    assign n1197 = n1092 ? n1133 : \pin_mux[11].pin_control [1];   // gpio_mux.v(78)
    assign n1198 = n1092 ? n1134 : \pin_mux[11].pin_control [0];   // gpio_mux.v(78)
    assign n1199 = n1092 ? n1135 : \pin_mux[10].pin_control [1];   // gpio_mux.v(78)
    assign n1200 = n1092 ? n1136 : \pin_mux[10].pin_control [0];   // gpio_mux.v(78)
    assign n1201 = n1092 ? n1137 : \pin_mux[9].pin_control [1];   // gpio_mux.v(78)
    assign n1202 = n1092 ? n1138 : \pin_mux[9].pin_control [0];   // gpio_mux.v(78)
    assign n1203 = n1092 ? n1139 : \pin_mux[8].pin_control [1];   // gpio_mux.v(78)
    assign n1204 = n1092 ? n1140 : \pin_mux[8].pin_control [0];   // gpio_mux.v(78)
    assign n1205 = n1092 ? n1141 : \pin_mux[7].pin_control [1];   // gpio_mux.v(78)
    assign n1206 = n1092 ? n1142 : \pin_mux[7].pin_control [0];   // gpio_mux.v(78)
    assign n1207 = n1092 ? n1143 : \pin_mux[6].pin_control [1];   // gpio_mux.v(78)
    assign n1208 = n1092 ? n1144 : \pin_mux[6].pin_control [0];   // gpio_mux.v(78)
    assign n1209 = n1092 ? n1145 : \pin_mux[5].pin_control [1];   // gpio_mux.v(78)
    assign n1210 = n1092 ? n1146 : \pin_mux[5].pin_control [0];   // gpio_mux.v(78)
    assign n1211 = n1092 ? n1147 : \pin_mux[4].pin_control [1];   // gpio_mux.v(78)
    assign n1212 = n1092 ? n1148 : \pin_mux[4].pin_control [0];   // gpio_mux.v(78)
    assign n1213 = n1092 ? n1149 : \pin_mux[3].pin_control [1];   // gpio_mux.v(78)
    assign n1214 = n1092 ? n1150 : \pin_mux[3].pin_control [0];   // gpio_mux.v(78)
    assign n1215 = n1092 ? n1151 : \pin_mux[2].pin_control [1];   // gpio_mux.v(78)
    assign n1216 = n1092 ? n1152 : \pin_mux[2].pin_control [0];   // gpio_mux.v(78)
    assign n1217 = n1092 ? n1153 : \pin_mux[1].pin_control [1];   // gpio_mux.v(78)
    assign n1218 = n1092 ? n1154 : \pin_mux[1].pin_control [0];   // gpio_mux.v(78)
    assign n1219 = n1092 ? n1155 : \pin_mux[0].pin_control [1];   // gpio_mux.v(78)
    assign n1220 = n1092 ? n1156 : \pin_mux[0].pin_control [0];   // gpio_mux.v(78)
    assign n1221 = sys_w ? n1157 : \pin_mux[31].pin_control [1];   // gpio_mux.v(77)
    assign n1222 = sys_w ? n1158 : \pin_mux[31].pin_control [0];   // gpio_mux.v(77)
    assign n1223 = sys_w ? n1159 : \pin_mux[30].pin_control [1];   // gpio_mux.v(77)
    assign n1224 = sys_w ? n1160 : \pin_mux[30].pin_control [0];   // gpio_mux.v(77)
    assign n1225 = sys_w ? n1161 : \pin_mux[29].pin_control [1];   // gpio_mux.v(77)
    assign n1226 = sys_w ? n1162 : \pin_mux[29].pin_control [0];   // gpio_mux.v(77)
    assign n1227 = sys_w ? n1163 : \pin_mux[28].pin_control [1];   // gpio_mux.v(77)
    assign n1228 = sys_w ? n1164 : \pin_mux[28].pin_control [0];   // gpio_mux.v(77)
    assign n1229 = sys_w ? n1165 : \pin_mux[27].pin_control [1];   // gpio_mux.v(77)
    assign n1230 = sys_w ? n1166 : \pin_mux[27].pin_control [0];   // gpio_mux.v(77)
    assign n1231 = sys_w ? n1167 : \pin_mux[26].pin_control [1];   // gpio_mux.v(77)
    assign n1232 = sys_w ? n1168 : \pin_mux[26].pin_control [0];   // gpio_mux.v(77)
    assign n1233 = sys_w ? n1169 : \pin_mux[25].pin_control [1];   // gpio_mux.v(77)
    assign n1234 = sys_w ? n1170 : \pin_mux[25].pin_control [0];   // gpio_mux.v(77)
    assign n1235 = sys_w ? n1171 : \pin_mux[24].pin_control [1];   // gpio_mux.v(77)
    assign n1236 = sys_w ? n1172 : \pin_mux[24].pin_control [0];   // gpio_mux.v(77)
    assign n1237 = sys_w ? n1173 : \pin_mux[23].pin_control [1];   // gpio_mux.v(77)
    assign n1238 = sys_w ? n1174 : \pin_mux[23].pin_control [0];   // gpio_mux.v(77)
    assign n1239 = sys_w ? n1175 : \pin_mux[22].pin_control [1];   // gpio_mux.v(77)
    assign n1240 = sys_w ? n1176 : \pin_mux[22].pin_control [0];   // gpio_mux.v(77)
    assign n1241 = sys_w ? n1177 : \pin_mux[21].pin_control [1];   // gpio_mux.v(77)
    assign n1242 = sys_w ? n1178 : \pin_mux[21].pin_control [0];   // gpio_mux.v(77)
    assign n1243 = sys_w ? n1179 : \pin_mux[20].pin_control [1];   // gpio_mux.v(77)
    assign n1244 = sys_w ? n1180 : \pin_mux[20].pin_control [0];   // gpio_mux.v(77)
    assign n1245 = sys_w ? n1181 : \pin_mux[19].pin_control [1];   // gpio_mux.v(77)
    assign n1246 = sys_w ? n1182 : \pin_mux[19].pin_control [0];   // gpio_mux.v(77)
    assign n1247 = sys_w ? n1183 : \pin_mux[18].pin_control [1];   // gpio_mux.v(77)
    assign n1248 = sys_w ? n1184 : \pin_mux[18].pin_control [0];   // gpio_mux.v(77)
    assign n1249 = sys_w ? n1185 : \pin_mux[17].pin_control [1];   // gpio_mux.v(77)
    assign n1250 = sys_w ? n1186 : \pin_mux[17].pin_control [0];   // gpio_mux.v(77)
    assign n1251 = sys_w ? n1187 : \pin_mux[16].pin_control [1];   // gpio_mux.v(77)
    assign n1252 = sys_w ? n1188 : \pin_mux[16].pin_control [0];   // gpio_mux.v(77)
    assign n1253 = sys_w ? n1189 : \pin_mux[15].pin_control [1];   // gpio_mux.v(77)
    assign n1254 = sys_w ? n1190 : \pin_mux[15].pin_control [0];   // gpio_mux.v(77)
    assign n1255 = sys_w ? n1191 : \pin_mux[14].pin_control [1];   // gpio_mux.v(77)
    assign n1256 = sys_w ? n1192 : \pin_mux[14].pin_control [0];   // gpio_mux.v(77)
    assign n1257 = sys_w ? n1193 : \pin_mux[13].pin_control [1];   // gpio_mux.v(77)
    assign n1258 = sys_w ? n1194 : \pin_mux[13].pin_control [0];   // gpio_mux.v(77)
    assign n1259 = sys_w ? n1195 : \pin_mux[12].pin_control [1];   // gpio_mux.v(77)
    assign n1260 = sys_w ? n1196 : \pin_mux[12].pin_control [0];   // gpio_mux.v(77)
    assign n1261 = sys_w ? n1197 : \pin_mux[11].pin_control [1];   // gpio_mux.v(77)
    assign n1262 = sys_w ? n1198 : \pin_mux[11].pin_control [0];   // gpio_mux.v(77)
    assign n1263 = sys_w ? n1199 : \pin_mux[10].pin_control [1];   // gpio_mux.v(77)
    assign n1264 = sys_w ? n1200 : \pin_mux[10].pin_control [0];   // gpio_mux.v(77)
    assign n1265 = sys_w ? n1201 : \pin_mux[9].pin_control [1];   // gpio_mux.v(77)
    assign n1266 = sys_w ? n1202 : \pin_mux[9].pin_control [0];   // gpio_mux.v(77)
    assign n1267 = sys_w ? n1203 : \pin_mux[8].pin_control [1];   // gpio_mux.v(77)
    assign n1268 = sys_w ? n1204 : \pin_mux[8].pin_control [0];   // gpio_mux.v(77)
    assign n1269 = sys_w ? n1205 : \pin_mux[7].pin_control [1];   // gpio_mux.v(77)
    assign n1270 = sys_w ? n1206 : \pin_mux[7].pin_control [0];   // gpio_mux.v(77)
    assign n1271 = sys_w ? n1207 : \pin_mux[6].pin_control [1];   // gpio_mux.v(77)
    assign n1272 = sys_w ? n1208 : \pin_mux[6].pin_control [0];   // gpio_mux.v(77)
    assign n1273 = sys_w ? n1209 : \pin_mux[5].pin_control [1];   // gpio_mux.v(77)
    assign n1274 = sys_w ? n1210 : \pin_mux[5].pin_control [0];   // gpio_mux.v(77)
    assign n1275 = sys_w ? n1211 : \pin_mux[4].pin_control [1];   // gpio_mux.v(77)
    assign n1276 = sys_w ? n1212 : \pin_mux[4].pin_control [0];   // gpio_mux.v(77)
    assign n1277 = sys_w ? n1213 : \pin_mux[3].pin_control [1];   // gpio_mux.v(77)
    assign n1278 = sys_w ? n1214 : \pin_mux[3].pin_control [0];   // gpio_mux.v(77)
    assign n1279 = sys_w ? n1215 : \pin_mux[2].pin_control [1];   // gpio_mux.v(77)
    assign n1280 = sys_w ? n1216 : \pin_mux[2].pin_control [0];   // gpio_mux.v(77)
    assign n1281 = sys_w ? n1217 : \pin_mux[1].pin_control [1];   // gpio_mux.v(77)
    assign n1282 = sys_w ? n1218 : \pin_mux[1].pin_control [0];   // gpio_mux.v(77)
    assign n1283 = sys_w ? n1219 : \pin_mux[0].pin_control [1];   // gpio_mux.v(77)
    assign n1284 = sys_w ? n1220 : \pin_mux[0].pin_control [0];   // gpio_mux.v(77)
    VERIFIC_DFFRS i1286 (.d(n1222), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[31].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1287 (.d(n1223), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[30].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1288 (.d(n1224), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[30].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1289 (.d(n1225), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[29].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1290 (.d(n1226), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[29].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1291 (.d(n1227), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[28].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1292 (.d(n1228), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[28].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1293 (.d(n1229), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[27].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1294 (.d(n1230), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[27].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1295 (.d(n1231), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[26].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1296 (.d(n1232), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[26].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1297 (.d(n1233), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[25].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1298 (.d(n1234), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[25].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1299 (.d(n1235), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[24].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1300 (.d(n1236), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[24].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1301 (.d(n1237), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[23].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1302 (.d(n1238), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[23].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1303 (.d(n1239), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[22].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1304 (.d(n1240), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[22].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1305 (.d(n1241), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[21].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1306 (.d(n1242), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[21].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1307 (.d(n1243), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[20].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1308 (.d(n1244), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[20].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1309 (.d(n1245), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[19].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1310 (.d(n1246), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[19].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1311 (.d(n1247), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[18].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1312 (.d(n1248), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[18].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1313 (.d(n1249), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[17].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1314 (.d(n1250), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[17].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1315 (.d(n1251), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[16].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1316 (.d(n1252), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[16].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1317 (.d(n1253), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[15].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1318 (.d(n1254), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[15].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1319 (.d(n1255), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[14].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1320 (.d(n1256), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[14].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1321 (.d(n1257), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[13].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1322 (.d(n1258), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[13].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1323 (.d(n1259), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[12].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1324 (.d(n1260), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[12].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1325 (.d(n1261), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[11].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1326 (.d(n1262), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[11].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1327 (.d(n1263), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[10].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1328 (.d(n1264), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[10].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1329 (.d(n1265), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[9].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1330 (.d(n1266), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[9].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1331 (.d(n1267), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[8].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1332 (.d(n1268), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[8].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1333 (.d(n1269), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[7].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1334 (.d(n1270), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[7].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1335 (.d(n1271), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[6].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1336 (.d(n1272), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[6].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1337 (.d(n1273), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[5].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1338 (.d(n1274), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[5].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1339 (.d(n1275), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[4].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1340 (.d(n1276), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[4].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1341 (.d(n1277), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[3].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1342 (.d(n1278), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[3].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1343 (.d(n1279), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[2].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1344 (.d(n1280), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[2].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1345 (.d(n1281), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[1].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1346 (.d(n1282), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[1].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1347 (.d(n1283), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[0].pin_control [1]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1348 (.d(n1284), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[0].pin_control [0]));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1349 (.d(n1424), .clk(clk), .s(1'b0), .r(1'b0), .q(n1349));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1350 (.d(n1438), .clk(clk), .s(1'b0), .r(1'b0), .q(n1350));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1351 (.d(n1452), .clk(clk), .s(1'b0), .r(1'b0), .q(n1351));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1352 (.d(n1466), .clk(clk), .s(1'b0), .r(1'b0), .q(n1352));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1353 (.d(n1480), .clk(clk), .s(1'b0), .r(1'b0), .q(n1353));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1354 (.d(n1494), .clk(clk), .s(1'b0), .r(1'b0), .q(n1354));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1355 (.d(n1508), .clk(clk), .s(1'b0), .r(1'b0), .q(n1355));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1356 (.d(n1522), .clk(clk), .s(1'b0), .r(1'b0), .q(n1356));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1357 (.d(n1536), .clk(clk), .s(1'b0), .r(1'b0), .q(n1357));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1358 (.d(n1550), .clk(clk), .s(1'b0), .r(1'b0), .q(n1358));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1359 (.d(n1564), .clk(clk), .s(1'b0), .r(1'b0), .q(n1359));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1360 (.d(n1578), .clk(clk), .s(1'b0), .r(1'b0), .q(n1360));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1361 (.d(n1592), .clk(clk), .s(1'b0), .r(1'b0), .q(n1361));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1362 (.d(n1606), .clk(clk), .s(1'b0), .r(1'b0), .q(n1362));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1363 (.d(n1620), .clk(clk), .s(1'b0), .r(1'b0), .q(n1363));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1364 (.d(n1634), .clk(clk), .s(1'b0), .r(1'b0), .q(n1364));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1365 (.d(n1648), .clk(clk), .s(1'b0), .r(1'b0), .q(n1365));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1366 (.d(n1662), .clk(clk), .s(1'b0), .r(1'b0), .q(n1366));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1367 (.d(n1676), .clk(clk), .s(1'b0), .r(1'b0), .q(n1367));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1368 (.d(n1690), .clk(clk), .s(1'b0), .r(1'b0), .q(n1368));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1369 (.d(n1704), .clk(clk), .s(1'b0), .r(1'b0), .q(n1369));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1370 (.d(n1718), .clk(clk), .s(1'b0), .r(1'b0), .q(n1370));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1371 (.d(n1732), .clk(clk), .s(1'b0), .r(1'b0), .q(n1371));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1372 (.d(n1746), .clk(clk), .s(1'b0), .r(1'b0), .q(n1372));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1373 (.d(n1760), .clk(clk), .s(1'b0), .r(1'b0), .q(n1373));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1374 (.d(n1774), .clk(clk), .s(1'b0), .r(1'b0), .q(n1374));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1375 (.d(n1788), .clk(clk), .s(1'b0), .r(1'b0), .q(n1375));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1376 (.d(n1802), .clk(clk), .s(1'b0), .r(1'b0), .q(n1376));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1377 (.d(n1816), .clk(clk), .s(1'b0), .r(1'b0), .q(n1377));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1378 (.d(n1830), .clk(clk), .s(1'b0), .r(1'b0), .q(n1378));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1379 (.d(n1844), .clk(clk), .s(1'b0), .r(1'b0), .q(n1379));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1380 (.d(n1858), .clk(clk), .s(1'b0), .r(1'b0), .q(n1380));   // gpio_mux.v(63)
    VERIFIC_DFFRS i1423 (.d(n1425), .clk(clk), .s(1'b0), .r(1'b0), .q(n1423));   // gpio_mux.v(63)
    not (n1416, rst) ;   // gpio_mux.v(63)
    and (n1421, sys_r, n964) ;   // gpio_mux.v(74)
    VERIFIC_DFFRS i1437 (.d(n1439), .clk(clk), .s(1'b0), .r(1'b0), .q(n1437));   // gpio_mux.v(63)
    assign n1424 = n1416 ? n965 : n1349;   // gpio_mux.v(63)
    assign n1425 = n1416 ? n1421 : n1423;   // gpio_mux.v(63)
    assign sys_r_line[31] = n1423 ? n1349 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1451 (.d(n1453), .clk(clk), .s(1'b0), .r(1'b0), .q(n1451));   // gpio_mux.v(63)
    assign n1438 = n1416 ? n966 : n1350;   // gpio_mux.v(63)
    assign n1439 = n1416 ? n1421 : n1437;   // gpio_mux.v(63)
    assign sys_r_line[30] = n1437 ? n1350 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1465 (.d(n1467), .clk(clk), .s(1'b0), .r(1'b0), .q(n1465));   // gpio_mux.v(63)
    assign n1452 = n1416 ? n967 : n1351;   // gpio_mux.v(63)
    assign n1453 = n1416 ? n1421 : n1451;   // gpio_mux.v(63)
    assign sys_r_line[29] = n1451 ? n1351 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1479 (.d(n1481), .clk(clk), .s(1'b0), .r(1'b0), .q(n1479));   // gpio_mux.v(63)
    assign n1466 = n1416 ? n968 : n1352;   // gpio_mux.v(63)
    assign n1467 = n1416 ? n1421 : n1465;   // gpio_mux.v(63)
    assign sys_r_line[28] = n1465 ? n1352 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1493 (.d(n1495), .clk(clk), .s(1'b0), .r(1'b0), .q(n1493));   // gpio_mux.v(63)
    assign n1480 = n1416 ? n969 : n1353;   // gpio_mux.v(63)
    assign n1481 = n1416 ? n1421 : n1479;   // gpio_mux.v(63)
    assign sys_r_line[27] = n1479 ? n1353 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1507 (.d(n1509), .clk(clk), .s(1'b0), .r(1'b0), .q(n1507));   // gpio_mux.v(63)
    assign n1494 = n1416 ? n970 : n1354;   // gpio_mux.v(63)
    assign n1495 = n1416 ? n1421 : n1493;   // gpio_mux.v(63)
    assign sys_r_line[26] = n1493 ? n1354 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1521 (.d(n1523), .clk(clk), .s(1'b0), .r(1'b0), .q(n1521));   // gpio_mux.v(63)
    assign n1508 = n1416 ? n971 : n1355;   // gpio_mux.v(63)
    assign n1509 = n1416 ? n1421 : n1507;   // gpio_mux.v(63)
    assign sys_r_line[25] = n1507 ? n1355 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1535 (.d(n1537), .clk(clk), .s(1'b0), .r(1'b0), .q(n1535));   // gpio_mux.v(63)
    assign n1522 = n1416 ? n972 : n1356;   // gpio_mux.v(63)
    assign n1523 = n1416 ? n1421 : n1521;   // gpio_mux.v(63)
    assign sys_r_line[24] = n1521 ? n1356 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1549 (.d(n1551), .clk(clk), .s(1'b0), .r(1'b0), .q(n1549));   // gpio_mux.v(63)
    assign n1536 = n1416 ? n973 : n1357;   // gpio_mux.v(63)
    assign n1537 = n1416 ? n1421 : n1535;   // gpio_mux.v(63)
    assign sys_r_line[23] = n1535 ? n1357 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1563 (.d(n1565), .clk(clk), .s(1'b0), .r(1'b0), .q(n1563));   // gpio_mux.v(63)
    assign n1550 = n1416 ? n974 : n1358;   // gpio_mux.v(63)
    assign n1551 = n1416 ? n1421 : n1549;   // gpio_mux.v(63)
    assign sys_r_line[22] = n1549 ? n1358 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1577 (.d(n1579), .clk(clk), .s(1'b0), .r(1'b0), .q(n1577));   // gpio_mux.v(63)
    assign n1564 = n1416 ? n975 : n1359;   // gpio_mux.v(63)
    assign n1565 = n1416 ? n1421 : n1563;   // gpio_mux.v(63)
    assign sys_r_line[21] = n1563 ? n1359 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1591 (.d(n1593), .clk(clk), .s(1'b0), .r(1'b0), .q(n1591));   // gpio_mux.v(63)
    assign n1578 = n1416 ? n976 : n1360;   // gpio_mux.v(63)
    assign n1579 = n1416 ? n1421 : n1577;   // gpio_mux.v(63)
    assign sys_r_line[20] = n1577 ? n1360 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1605 (.d(n1607), .clk(clk), .s(1'b0), .r(1'b0), .q(n1605));   // gpio_mux.v(63)
    assign n1592 = n1416 ? n977 : n1361;   // gpio_mux.v(63)
    assign n1593 = n1416 ? n1421 : n1591;   // gpio_mux.v(63)
    assign sys_r_line[19] = n1591 ? n1361 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1619 (.d(n1621), .clk(clk), .s(1'b0), .r(1'b0), .q(n1619));   // gpio_mux.v(63)
    assign n1606 = n1416 ? n978 : n1362;   // gpio_mux.v(63)
    assign n1607 = n1416 ? n1421 : n1605;   // gpio_mux.v(63)
    assign sys_r_line[18] = n1605 ? n1362 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1633 (.d(n1635), .clk(clk), .s(1'b0), .r(1'b0), .q(n1633));   // gpio_mux.v(63)
    assign n1620 = n1416 ? n979 : n1363;   // gpio_mux.v(63)
    assign n1621 = n1416 ? n1421 : n1619;   // gpio_mux.v(63)
    assign sys_r_line[17] = n1619 ? n1363 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1647 (.d(n1649), .clk(clk), .s(1'b0), .r(1'b0), .q(n1647));   // gpio_mux.v(63)
    assign n1634 = n1416 ? n980 : n1364;   // gpio_mux.v(63)
    assign n1635 = n1416 ? n1421 : n1633;   // gpio_mux.v(63)
    assign sys_r_line[16] = n1633 ? n1364 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1661 (.d(n1663), .clk(clk), .s(1'b0), .r(1'b0), .q(n1661));   // gpio_mux.v(63)
    assign n1648 = n1416 ? n981 : n1365;   // gpio_mux.v(63)
    assign n1649 = n1416 ? n1421 : n1647;   // gpio_mux.v(63)
    assign sys_r_line[15] = n1647 ? n1365 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1675 (.d(n1677), .clk(clk), .s(1'b0), .r(1'b0), .q(n1675));   // gpio_mux.v(63)
    assign n1662 = n1416 ? n982 : n1366;   // gpio_mux.v(63)
    assign n1663 = n1416 ? n1421 : n1661;   // gpio_mux.v(63)
    assign sys_r_line[14] = n1661 ? n1366 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1689 (.d(n1691), .clk(clk), .s(1'b0), .r(1'b0), .q(n1689));   // gpio_mux.v(63)
    assign n1676 = n1416 ? n983 : n1367;   // gpio_mux.v(63)
    assign n1677 = n1416 ? n1421 : n1675;   // gpio_mux.v(63)
    assign sys_r_line[13] = n1675 ? n1367 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1703 (.d(n1705), .clk(clk), .s(1'b0), .r(1'b0), .q(n1703));   // gpio_mux.v(63)
    assign n1690 = n1416 ? n984 : n1368;   // gpio_mux.v(63)
    assign n1691 = n1416 ? n1421 : n1689;   // gpio_mux.v(63)
    assign sys_r_line[12] = n1689 ? n1368 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1717 (.d(n1719), .clk(clk), .s(1'b0), .r(1'b0), .q(n1717));   // gpio_mux.v(63)
    assign n1704 = n1416 ? n985 : n1369;   // gpio_mux.v(63)
    assign n1705 = n1416 ? n1421 : n1703;   // gpio_mux.v(63)
    assign sys_r_line[11] = n1703 ? n1369 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1731 (.d(n1733), .clk(clk), .s(1'b0), .r(1'b0), .q(n1731));   // gpio_mux.v(63)
    assign n1718 = n1416 ? n986 : n1370;   // gpio_mux.v(63)
    assign n1719 = n1416 ? n1421 : n1717;   // gpio_mux.v(63)
    assign sys_r_line[10] = n1717 ? n1370 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1745 (.d(n1747), .clk(clk), .s(1'b0), .r(1'b0), .q(n1745));   // gpio_mux.v(63)
    assign n1732 = n1416 ? n987 : n1371;   // gpio_mux.v(63)
    assign n1733 = n1416 ? n1421 : n1731;   // gpio_mux.v(63)
    assign sys_r_line[9] = n1731 ? n1371 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1759 (.d(n1761), .clk(clk), .s(1'b0), .r(1'b0), .q(n1759));   // gpio_mux.v(63)
    assign n1746 = n1416 ? n988 : n1372;   // gpio_mux.v(63)
    assign n1747 = n1416 ? n1421 : n1745;   // gpio_mux.v(63)
    assign sys_r_line[8] = n1745 ? n1372 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1773 (.d(n1775), .clk(clk), .s(1'b0), .r(1'b0), .q(n1773));   // gpio_mux.v(63)
    assign n1760 = n1416 ? n989 : n1373;   // gpio_mux.v(63)
    assign n1761 = n1416 ? n1421 : n1759;   // gpio_mux.v(63)
    assign sys_r_line[7] = n1759 ? n1373 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1787 (.d(n1789), .clk(clk), .s(1'b0), .r(1'b0), .q(n1787));   // gpio_mux.v(63)
    assign n1774 = n1416 ? n990 : n1374;   // gpio_mux.v(63)
    assign n1775 = n1416 ? n1421 : n1773;   // gpio_mux.v(63)
    assign sys_r_line[6] = n1773 ? n1374 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1801 (.d(n1803), .clk(clk), .s(1'b0), .r(1'b0), .q(n1801));   // gpio_mux.v(63)
    assign n1788 = n1416 ? n991 : n1375;   // gpio_mux.v(63)
    assign n1789 = n1416 ? n1421 : n1787;   // gpio_mux.v(63)
    assign sys_r_line[5] = n1787 ? n1375 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1815 (.d(n1817), .clk(clk), .s(1'b0), .r(1'b0), .q(n1815));   // gpio_mux.v(63)
    assign n1802 = n1416 ? n992 : n1376;   // gpio_mux.v(63)
    assign n1803 = n1416 ? n1421 : n1801;   // gpio_mux.v(63)
    assign sys_r_line[4] = n1801 ? n1376 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1829 (.d(n1831), .clk(clk), .s(1'b0), .r(1'b0), .q(n1829));   // gpio_mux.v(63)
    assign n1816 = n1416 ? n993 : n1377;   // gpio_mux.v(63)
    assign n1817 = n1416 ? n1421 : n1815;   // gpio_mux.v(63)
    assign sys_r_line[3] = n1815 ? n1377 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1843 (.d(n1845), .clk(clk), .s(1'b0), .r(1'b0), .q(n1843));   // gpio_mux.v(63)
    assign n1830 = n1416 ? n994 : n1378;   // gpio_mux.v(63)
    assign n1831 = n1416 ? n1421 : n1829;   // gpio_mux.v(63)
    assign sys_r_line[2] = n1829 ? n1378 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1857 (.d(n1859), .clk(clk), .s(1'b0), .r(1'b0), .q(n1857));   // gpio_mux.v(63)
    assign n1844 = n1416 ? n995 : n1379;   // gpio_mux.v(63)
    assign n1845 = n1416 ? n1421 : n1843;   // gpio_mux.v(63)
    assign sys_r_line[1] = n1843 ? n1379 : 1'bz;   // gpio_mux.v(58)
    assign n1858 = n1416 ? n996 : n1380;   // gpio_mux.v(63)
    assign n1859 = n1416 ? n1421 : n1857;   // gpio_mux.v(63)
    assign sys_r_line[0] = n1857 ? n1380 : 1'bz;   // gpio_mux.v(58)
    VERIFIC_DFFRS i1285 (.d(n1221), .clk(clk), .s(1'b0), .r(rst), .q(\pin_mux[31].pin_control [1]));   // gpio_mux.v(63)
    
endmodule
