
//
// Verific Verilog Description of module test_pipeline_assembly
//

module test_pipeline_assembly (ram_w_addr, ram_r_addr, ram_w_line, ram_read, 
            ram_write, sys_w_addr, sys_r_addr, sys_w_line, sys_read, 
            sys_write, lr, sp, pc, st, word, ram_r_line, sys_r_line, 
            clk, rst);   // test_pipeline_assembly.v(32)
    output [31:0]ram_w_addr;   // test_pipeline_assembly.v(37)
    output [31:0]ram_r_addr;   // test_pipeline_assembly.v(37)
    output [31:0]ram_w_line;   // test_pipeline_assembly.v(38)
    output ram_read;   // test_pipeline_assembly.v(40)
    output ram_write;   // test_pipeline_assembly.v(40)
    output [31:0]sys_w_addr;   // test_pipeline_assembly.v(42)
    output [31:0]sys_r_addr;   // test_pipeline_assembly.v(42)
    output [31:0]sys_w_line;   // test_pipeline_assembly.v(43)
    output sys_read;   // test_pipeline_assembly.v(45)
    output sys_write;   // test_pipeline_assembly.v(45)
    output [31:0]lr;   // test_pipeline_assembly.v(47)
    output [31:0]sp;   // test_pipeline_assembly.v(47)
    output [31:0]pc;   // test_pipeline_assembly.v(47)
    output [31:0]st;   // test_pipeline_assembly.v(47)
    input [31:0]word;   // test_pipeline_assembly.v(33)
    input [31:0]ram_r_line;   // test_pipeline_assembly.v(39)
    input [31:0]sys_r_line;   // test_pipeline_assembly.v(44)
    input clk;   // test_pipeline_assembly.v(35)
    input rst;   // test_pipeline_assembly.v(35)
    
    wire [31:0]reg_c;   // test_pipeline_assembly.v(54)
    wire [31:0]reg_d;   // test_pipeline_assembly.v(54)
    wire [4:0]reg_a_a;   // test_pipeline_assembly.v(55)
    wire [4:0]reg_a_b;   // test_pipeline_assembly.v(55)
    wire [4:0]reg_a_c;   // test_pipeline_assembly.v(55)
    wire [4:0]reg_a_d;   // test_pipeline_assembly.v(55)
    wire [1:0]reg_read;   // test_pipeline_assembly.v(56)
    wire [1:0]reg_write;   // test_pipeline_assembly.v(56)
    wire [31:0]reg_stin;   // test_pipeline_assembly.v(59)
    wire reg_stwr;   // test_pipeline_assembly.v(60)
    wire reg_pcincr;   // test_pipeline_assembly.v(61)
    wire [31:0]e_a;   // test_pipeline_assembly.v(65)
    wire [31:0]e_b;   // test_pipeline_assembly.v(65)
    wire [7:0]e_alu_op;   // test_pipeline_assembly.v(66)
    wire [3:0]e_cond;   // test_pipeline_assembly.v(67)
    wire [3:0]e_write_flags;   // test_pipeline_assembly.v(68)
    wire e_swp;   // test_pipeline_assembly.v(69)
    wire e_is_cond;   // test_pipeline_assembly.v(70)
    wire [31:0]m_a1;   // test_pipeline_assembly.v(72)
    wire [31:0]m_a2;   // test_pipeline_assembly.v(72)
    wire [3:0]m_r1_op;   // test_pipeline_assembly.v(73)
    wire [3:0]m_r2_op;   // test_pipeline_assembly.v(73)
    wire [4:0]r_a1;   // test_pipeline_assembly.v(75)
    wire [4:0]r_a2;   // test_pipeline_assembly.v(75)
    wire [3:0]r_op;   // test_pipeline_assembly.v(76)
    wire d_pass;   // test_pipeline_assembly.v(78)
    wire d_pcincr;   // test_pipeline_assembly.v(79)
    wire [31:0]d_r1;   // test_pipeline_assembly.v(87)
    wire [31:0]d_r2;   // test_pipeline_assembly.v(87)
    wire d_hazard;   // test_pipeline_assembly.v(88)
    wire [31:0]pi_m_a1;   // test_pipeline_assembly.v(99)
    wire [31:0]pi_m_a2;   // test_pipeline_assembly.v(99)
    wire [3:0]pi_m_r1_op;   // test_pipeline_assembly.v(100)
    wire [3:0]pi_m_r2_op;   // test_pipeline_assembly.v(100)
    wire [4:0]pi_r_a1;   // test_pipeline_assembly.v(102)
    wire [4:0]pi_r_a2;   // test_pipeline_assembly.v(102)
    wire [3:0]pi_r_op;   // test_pipeline_assembly.v(103)
    wire [31:0]ex_a;   // test_pipeline_assembly.v(113)
    wire [31:0]ex_b;   // test_pipeline_assembly.v(113)
    wire [7:0]ex_alu_op;   // test_pipeline_assembly.v(115)
    wire ex_is_cond;   // test_pipeline_assembly.v(116)
    wire [3:0]ex_cond;   // test_pipeline_assembly.v(117)
    wire [3:0]ex_write_flags;   // test_pipeline_assembly.v(118)
    wire ex_swp;   // test_pipeline_assembly.v(119)
    wire ex_cres;   // test_pipeline_assembly.v(124)
    wire sr_n;   // test_pipeline_assembly.v(128)
    wire sr_z;   // test_pipeline_assembly.v(128)
    wire sr_c;   // test_pipeline_assembly.v(128)
    wire sr_v;   // test_pipeline_assembly.v(128)
    wire sr_cc;   // test_pipeline_assembly.v(129)
    wire [4:0]ex_r_a1;   // test_pipeline_assembly.v(141)
    wire [4:0]ex_r_a2;   // test_pipeline_assembly.v(141)
    wire [3:0]ex_r_op;   // test_pipeline_assembly.v(142)
    wire [31:0]mop_r1;   // test_pipeline_assembly.v(146)
    wire [31:0]mop_r2;   // test_pipeline_assembly.v(146)
    wire [31:0]mop_a1;   // test_pipeline_assembly.v(147)
    wire [31:0]mop_a2;   // test_pipeline_assembly.v(147)
    wire [3:0]mop_r1_op;   // test_pipeline_assembly.v(149)
    wire [3:0]mop_r2_op;   // test_pipeline_assembly.v(149)
    wire [4:0]mop_r_a1;   // test_pipeline_assembly.v(169)
    wire [4:0]mop_r_a2;   // test_pipeline_assembly.v(169)
    wire [3:0]mop_r_op;   // test_pipeline_assembly.v(170)
    wire mop_proceed2;   // test_pipeline_assembly.v(171)
    wire [31:0]rwb_r1;   // test_pipeline_assembly.v(175)
    wire [31:0]rwb_r2;   // test_pipeline_assembly.v(175)
    wire ex_hazard;   // test_pipeline_assembly.v(190)
    wire mem_hazard;   // test_pipeline_assembly.v(192)
    
    reg32_2x2_pc rf0 (.rd0({d_r1}), .rd1({d_r2}), .ra0({reg_a_a}), .ra1({reg_a_b}), 
            .wa0({reg_a_c}), .wa1({reg_a_d}), .wd0({reg_c}), .wd1({reg_d}), 
            .read({reg_read}), .write({reg_write}), .clk(clk), .rst(rst), 
            .lrout({lr}), .spout({sp}), .stout({st}), .pcout({pc}), 
            .stin({reg_stin}), .stwr(reg_stwr), .pcincr(reg_pcincr));   // test_pipeline_assembly.v(62)
    insn_decoder dec0 (.e_a({e_a}), .e_b({e_b}), .e_alu_op({e_alu_op}), 
            .e_is_cond(e_is_cond), .e_cond({e_cond}), .e_write_flags({e_write_flags}), 
            .e_swp(e_swp), .m_a1({m_a1}), .m_a2({m_a2}), .m_r1_op({m_r1_op}), 
            .m_r2_op({m_r2_op}), .r_a1({r_a1}), .r_a2({r_a2}), .r_op({r_op}), 
            .d_pass(d_pass), .d_pcincr(d_pcincr), .r_r1_addr({reg_a_a}), 
            .r_r2_addr({reg_a_b}), .r_read({reg_read}), .word({word}), 
            .r1({d_r1}), .r2({d_r2}), .hazard(d_hazard), .rst(rst), 
            .clk(clk));   // test_pipeline_assembly.v(89)
    pipeline_interface pi0 (.qe_a({ex_a}), .qe_b({ex_b}), .qe_alu_op({ex_alu_op}), 
            .qe_is_cond(ex_is_cond), .qe_cond({ex_cond}), .qe_write_flags({ex_write_flags}), 
            .qe_swp(ex_swp), .qm_a1({pi_m_a1}), .qm_a2({pi_m_a2}), .qm_r1_op({pi_m_r1_op}), 
            .qm_r2_op({pi_m_r2_op}), .qr_a1({pi_r_a1}), .qr_a2({pi_r_a2}), 
            .qr_op({pi_r_op}), .qd_pcincr(reg_pcincr), .e_a({e_a}), .e_b({e_b}), 
            .e_alu_op({e_alu_op}), .e_is_cond(e_is_cond), .e_cond({e_cond}), 
            .e_write_flags({e_write_flags}), .e_swp(e_swp), .m_a1({m_a1}), 
            .m_a2({m_a2}), .m_r1_op({m_r1_op}), .m_r2_op({m_r2_op}), .r_a1({r_a1}), 
            .r_a2({r_a2}), .r_op({r_op}), .d_pass(d_pass), .d_pcincr(d_pcincr), 
            .clk(clk), .rst(rst));   // test_pipeline_assembly.v(108)
    execute ex0 (.r1({mop_r1}), .r2({mop_r2}), .cres(ex_cres), .n(sr_n), 
            .z(sr_z), .c(sr_c), .v(sr_v), .cc(sr_cc), .a({ex_a}), 
            .b({ex_b}), .alu_op({ex_alu_op}), .is_cond(ex_is_cond), .cond({ex_cond}), 
            .write_flags({ex_write_flags}), .st({st}), .swp(ex_swp), .clk(clk), 
            .rst(rst));   // test_pipeline_assembly.v(125)
    status_register_adaptor sr0 (.st({reg_stin}), .stwr(reg_stwr), .n(sr_n), 
            .z(sr_z), .c(sr_c), .v(sr_v), .cc(sr_cc));   // test_pipeline_assembly.v(135)
    execute_stage_passthrough exh0 (.qm_a1({mop_a1}), .qm_a2({mop_a2}), 
            .qm_r1_op({mop_r1_op}), .qm_r2_op({mop_r2_op}), .qr_a1({ex_r_a1}), 
            .qr_a2({ex_r_a2}), .qr_op({ex_r_op}), .m_a1({pi_m_a1}), .m_a2({pi_m_a2}), 
            .m_r1_op({pi_m_r1_op}), .m_r2_op({pi_m_r2_op}), .r_a1({pi_r_a1}), 
            .r_a2({pi_r_a2}), .r_op({pi_r_op}), .clk(clk), .rst(rst));   // test_pipeline_assembly.v(143)
    memory_op mop0 (.m1({rwb_r1}), .m2({rwb_r2}), .ram_w_addr({ram_w_addr}), 
            .ram_r_addr({ram_r_addr}), .ram_w(ram_write), .ram_r(ram_read), 
            .ram_w_line({ram_w_line}), .sys_w_addr({sys_w_addr}), .sys_r_addr({sys_r_addr}), 
            .sys_w(sys_write), .sys_r(sys_read), .sys_w_line({sys_w_line}), 
            .r1({mop_r1}), .r2({mop_r2}), .a1({mop_a1}), .a2({mop_a2}), 
            .r1_op({mop_r1_op}), .r2_op({mop_r2_op}), .ram_r_line({ram_r_line}), 
            .sys_r_line({sys_r_line}), .proceed(ex_cres), .clk(clk), .rst(rst));   // test_pipeline_assembly.v(167)
    memory_op_stage_passthrough moph0 (.q_a1({mop_r_a1}), .q_a2({mop_r_a2}), 
            .q_op({mop_r_op}), .q_proceed(mop_proceed2), .a1({ex_r_a1}), 
            .a2({ex_r_a2}), .op({ex_r_op}), .proceed(ex_cres), .clk(clk), 
            .rst(rst));   // test_pipeline_assembly.v(172)
    register_wb rwb0 (.write({reg_write}), .wr1({reg_c}), .wr2({reg_d}), 
            .wa1({reg_a_c}), .wa2({reg_a_d}), .r1({rwb_r1}), .r2({rwb_r2}), 
            .a1({mop_r_a1}), .a2({mop_r_a2}), .op({mop_r_op}), .proceed(mop_proceed2), 
            .clk(clk), .rst(rst));   // test_pipeline_assembly.v(188)
    reg_hazard_checker hz0 (.ex_hazard(ex_hazard), .mem_hazard(mem_hazard), 
            .ex_r1_a({ex_r_a1}), .ex_r2_a({ex_r_a2}), .ex_r_op({ex_r_op}), 
            .ex_proceed(ex_cres), .mem_r1_a({mop_r_a1}), .mem_r2_a({mop_r_a2}), 
            .mem_r_op({mop_r_op}), .mem_proceed(mop_proceed2), .reg_r1_a({reg_a_c}), 
            .reg_r2_a({reg_a_d}), .reg_write({reg_write}), .dec_r1_addr({reg_a_a}), 
            .dec_r2_addr({reg_a_b}), .dec_r_read({reg_read}));   // test_pipeline_assembly.v(193)
    or (d_hazard, ex_hazard, mem_hazard) ;   // test_pipeline_assembly.v(197)
    
endmodule

//
// Verific Verilog Description of module reg32_2x2_pc
//

module reg32_2x2_pc (rd0, rd1, ra0, ra1, wa0, wa1, wd0, wd1, 
            read, write, clk, rst, lrout, spout, stout, pcout, 
            stin, stwr, pcincr);   // regs.v(4)
    output [31:0]rd0;   // regs.v(17)
    output [31:0]rd1;   // regs.v(17)
    input [4:0]ra0;   // regs.v(8)
    input [4:0]ra1;   // regs.v(8)
    input [4:0]wa0;   // regs.v(9)
    input [4:0]wa1;   // regs.v(9)
    input [31:0]wd0;   // regs.v(11)
    input [31:0]wd1;   // regs.v(11)
    input [1:0]read;   // regs.v(13)
    input [1:0]write;   // regs.v(13)
    input clk;   // regs.v(15)
    input rst;   // regs.v(15)
    output [31:0]lrout;   // regs.v(21)
    output [31:0]spout;   // regs.v(21)
    output [31:0]stout;   // regs.v(21)
    output [31:0]pcout;   // regs.v(21)
    input [31:0]stin;   // regs.v(22)
    input stwr;   // regs.v(23)
    input pcincr;   // regs.v(23)
    
    wire [31:0]\regs[27] ;   // regs.v(19)
    wire [31:0]\regs[26] ;   // regs.v(19)
    wire [31:0]\regs[25] ;   // regs.v(19)
    wire [31:0]\regs[24] ;   // regs.v(19)
    wire [31:0]\regs[23] ;   // regs.v(19)
    wire [31:0]\regs[22] ;   // regs.v(19)
    wire [31:0]\regs[21] ;   // regs.v(19)
    wire [31:0]\regs[20] ;   // regs.v(19)
    wire [31:0]\regs[19] ;   // regs.v(19)
    wire [31:0]\regs[18] ;   // regs.v(19)
    wire [31:0]\regs[17] ;   // regs.v(19)
    wire [31:0]\regs[16] ;   // regs.v(19)
    wire [31:0]\regs[15] ;   // regs.v(19)
    wire [31:0]\regs[14] ;   // regs.v(19)
    wire [31:0]\regs[13] ;   // regs.v(19)
    wire [31:0]\regs[12] ;   // regs.v(19)
    wire [31:0]\regs[11] ;   // regs.v(19)
    wire [31:0]\regs[10] ;   // regs.v(19)
    wire [31:0]\regs[9] ;   // regs.v(19)
    wire [31:0]\regs[8] ;   // regs.v(19)
    wire [31:0]\regs[7] ;   // regs.v(19)
    wire [31:0]\regs[6] ;   // regs.v(19)
    wire [31:0]\regs[5] ;   // regs.v(19)
    wire [31:0]\regs[4] ;   // regs.v(19)
    wire [31:0]\regs[3] ;   // regs.v(19)
    wire [31:0]\regs[2] ;   // regs.v(19)
    wire [31:0]\regs[1] ;   // regs.v(19)
    wire [31:0]\regs[0] ;   // regs.v(19)
    
    wire n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
        n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
        n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, 
        n99, n100, n101, n102, n103, n104, n105, n106, n107, 
        n108, n109, n110, n111, n112, n113, n114, n115, n116, 
        n117, n118, n119, n120, n121, n122, n123, n124, n125, 
        n126, n127, n128, n129, n130, n131, n132, n133, n134, 
        n135, n136, n137, n138, n139, n140, n141, n142, n143, 
        n144, n145, n146, n147, n148, n149, n150, n151, n152, 
        n153, n154, n155, n156, n157, n158, n159, n160, n161, 
        n162, n163, n164, n165, n166, n167, n168, n169, n170, 
        n171, n172, n173, n174, n175, n176, n177, n178, n179, 
        n180, n181, n182, n183, n184, n185, n186, n187, n188, 
        n189, n190, n191, n192, n193, n194, n195, n196, n197, 
        n198, n199, n200, n201, n202, n203, n204, n205, n206, 
        n207, n208, n209, n210, n211, n212, n213, n214, n215, 
        n216, n217, n218, n219, n220, n221, n222, n223, n224, 
        n225, n226, n227, n228, n229, n230, n231, n232, n233, 
        n234, n235, n236, n237, n238, n239, n240, n241, n242, 
        n243, n244, n245, n246, n247, n248, n249, n250, n251, 
        n252, n253, n254, n255, n256, n257, n258, n259, n260, 
        n261, n262, n263, n264, n265, n266, n267, n268, n269, 
        n270, n271, n272, n273, n274, n275, n276, n277, n278, 
        n279, n280, n281, n282, n283, n284, n285, n286, n287, 
        n288, n289, n290, n291, n292, n293, n294, n295, n296, 
        n297, n298, n299, n300, n301, n302, n303, n304, n305, 
        n306, n307, n308, n309, n310, n311, n312, n313, n314, 
        n315, n316, n317, n318, n319, n320, n321, n322, n323, 
        n324, n325, n326, n327, n328, n329, n330, n331, n332, 
        n333, n334, n335, n336, n337, n338, n339, n340, n341, 
        n342, n343, n344, n345, n346, n347, n348, n349, n350, 
        n351, n352, n353, n354, n355, n356, n357, n358, n359, 
        n360, n361, n362, n363, n364, n365, n366, n367, n368, 
        n369, n370, n371, n372, n373, n374, n375, n376, n377, 
        n378, n379, n380, n381, n382, n383, n384, n385, n386, 
        n387, n388, n389, n390, n391, n392, n393, n394, n395, 
        n396, n397, n398, n399, n400, n401, n402, n403, n404, 
        n405, n406, n407, n408, n409, n410, n411, n412, n413, 
        n414, n415, n416, n417, n418, n419, n420, n421, n422, 
        n423, n424, n425, n426, n427, n428, n429, n430, n431, 
        n432, n433, n434, n435, n436, n437, n438, n439, n440, 
        n441, n442, n443, n444, n445, n446, n447, n448, n449, 
        n450, n451, n452, n453, n454, n455, n456, n457, n458, 
        n459, n460, n461, n462, n463, n464, n465, n466, n467, 
        n468, n469, n470, n471, n472, n473, n474, n475, n476, 
        n477, n478, n479, n480, n481, n482, n483, n484, n485, 
        n486, n487, n488, n489, n490, n491, n492, n493, n494, 
        n495, n496, n497, n498, n499, n500, n501, n502, n503, 
        n504, n505, n506, n507, n508, n509, n510, n511, n512, 
        n513, n514, n515, n516, n517, n518, n519, n520, n521, 
        n522, n523, n524, n525, n526, n527, n528, n529, n530, 
        n531, n532, n533, n534, n535, n536, n537, n538, n539, 
        n540, n541, n542, n543, n544, n545, n546, n547, n548, 
        n549, n550, n551, n552, n553, n554, n555, n556, n557, 
        n558, n559, n560, n561, n562, n563, n564, n565, n566, 
        n567, n568, n569, n570, n571, n572, n573, n574, n575, 
        n576, n577, n578, n579, n580, n581, n582, n583, n584, 
        n585, n586, n587, n588, n589, n590, n591, n592, n593, 
        n594, n595, n596, n597, n598, n599, n600, n601, n602, 
        n603, n604, n605, n606, n607, n608, n609, n610, n611, 
        n612, n613, n614, n615, n616, n617, n618, n619, n620, 
        n621, n622, n623, n624, n625, n626, n627, n628, n629, 
        n630, n631, n632, n633, n634, n635, n636, n637, n638, 
        n639, n640, n641, n642, n643, n644, n645, n646, n647, 
        n648, n649, n650, n651, n652, n653, n654, n655, n656, 
        n657, n658, n659, n660, n661, n662, n663, n664, n665, 
        n666, n667, n668, n669, n670, n671, n672, n673, n674, 
        n675, n676, n677, n678, n679, n680, n681, n682, n683, 
        n684, n685, n686, n687, n688, n689, n690, n691, n692, 
        n693, n694, n695, n696, n697, n698, n699, n700, n701, 
        n702, n703, n704, n705, n706, n707, n708, n709, n710, 
        n711, n712, n713, n714, n715, n716, n717, n718, n719, 
        n720, n721, n722, n723, n724, n725, n726, n727, n728, 
        n729, n730, n731, n732, n733, n734, n735, n736, n737, 
        n738, n739, n740, n741, n742, n743, n744, n745, n746, 
        n747, n748, n749, n750, n751, n752, n753, n754, n755, 
        n756, n757, n758, n759, n760, n761, n762, n763, n764, 
        n765, n766, n767, n768, n769, n770, n771, n772, n773, 
        n774, n775, n776, n777, n778, n779, n780, n781, n782, 
        n783, n784, n785, n786, n787, n788, n789, n790, n791, 
        n792, n793, n794, n795, n796, n797, n798, n799, n800, 
        n801, n802, n803, n804, n805, n806, n807, n808, n809, 
        n810, n811, n812, n813, n814, n815, n816, n817, n818, 
        n819, n820, n821, n822, n823, n824, n825, n826, n827, 
        n828, n829, n830, n831, n832, n833, n834, n835, n836, 
        n837, n838, n839, n840, n841, n842, n843, n844, n845, 
        n846, n847, n848, n849, n850, n851, n852, n853, n854, 
        n855, n856, n857, n858, n859, n860, n861, n862, n863, 
        n864, n865, n866, n867, n868, n869, n870, n871, n872, 
        n873, n874, n875, n876, n877, n878, n879, n880, n881, 
        n882, n883, n884, n885, n886, n887, n888, n889, n890, 
        n891, n892, n893, n894, n895, n896, n897, n898, n899, 
        n900, n901, n902, n903, n904, n905, n906, n907, n908, 
        n909, n910, n911, n912, n913, n914, n915, n916, n917, 
        n918, n919, n920, n921, n922, n923, n924, n925, n926, 
        n927, n928, n929, n930, n931, n932, n933, n934, n935, 
        n936, n937, n938, n939, n940, n941, n942, n943, n944, 
        n945, n946, n947, n948, n949, n950, n951, n952, n953, 
        n954, n955, n956, n957, n958, n959, n960, n961, n962, 
        n963, n964, n965, n966, n967, n968, n969, n970, n971, 
        n972, n973, n974, n975, n976, n977, n978, n979, n980, 
        n981, n982, n983, n984, n985, n986, n987, n988, n989, 
        n990, n991, n992, n993, n994, n995, n996, n997, n998, 
        n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, 
        n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, 
        n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
        n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
        n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, 
        n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, 
        n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, 
        n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
        n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, 
        n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, 
        n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, 
        n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, 
        n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
        n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, 
        n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, 
        n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, 
        n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, 
        n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
        n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, 
        n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, 
        n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
        n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, 
        n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
        n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, 
        n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, 
        n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
        n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, 
        n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
        n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, 
        n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, 
        n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
        n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, 
        n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
        n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, 
        n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, 
        n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
        n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, 
        n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
        n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, 
        n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, 
        n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
        n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, 
        n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
        n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, 
        n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, 
        n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
        n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, 
        n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, 
        n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, 
        n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, 
        n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
        n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, 
        n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, 
        n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, 
        n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, 
        n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
        n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, 
        n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, 
        n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, 
        n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, 
        n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
        n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, 
        n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
        n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, 
        n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, 
        n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
        n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, 
        n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
        n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, 
        n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, 
        n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
        n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, 
        n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
        n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, 
        n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, 
        n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
        n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, 
        n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
        n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, 
        n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, 
        n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
        n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, 
        n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, 
        n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, 
        n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, 
        n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
        n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, 
        n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, 
        n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, 
        n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, 
        n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
        n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, 
        n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, 
        n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, 
        n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, 
        n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
        n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, 
        n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, 
        n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, 
        n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, 
        n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
        n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, 
        n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
        n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, 
        n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, 
        n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
        n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, 
        n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
        n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, 
        n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, 
        n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
        n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, 
        n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, 
        n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, 
        n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, 
        n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
        n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, 
        n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, 
        n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, 
        n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, 
        n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
        n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, 
        n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
        n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, 
        n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, 
        n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
        n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, 
        n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
        n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, 
        n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, 
        n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
        n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, 
        n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
        n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, 
        n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, 
        n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
        n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, 
        n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
        n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, 
        n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, 
        n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
        n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, 
        n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
        n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, 
        n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, 
        n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
        n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, 
        n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
        n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, 
        n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, 
        n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, 
        n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, 
        n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
        n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, 
        n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, 
        n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, 
        n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, 
        n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
        n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, 
        n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, 
        n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, 
        n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, 
        n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, 
        n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, 
        n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, 
        n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, 
        n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, 
        n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, 
        n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, 
        n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, 
        n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, 
        n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, 
        n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, 
        n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, 
        n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, 
        n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, 
        n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, 
        n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
        n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, 
        n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, 
        n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, 
        n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, 
        n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, 
        n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, 
        n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, 
        n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, 
        n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, 
        n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, 
        n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, 
        n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, 
        n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, 
        n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, 
        n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, 
        n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, 
        n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, 
        n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, 
        n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, 
        n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, 
        n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, 
        n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, 
        n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, 
        n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, 
        n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, 
        n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, 
        n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, 
        n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, 
        n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, 
        n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, 
        n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, 
        n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, 
        n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, 
        n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, 
        n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, 
        n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, 
        n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, 
        n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, 
        n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, 
        n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, 
        n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, 
        n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, 
        n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, 
        n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, 
        n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, 
        n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, 
        n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, 
        n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, 
        n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, 
        n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, 
        n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, 
        n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, 
        n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, 
        n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, 
        n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, 
        n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, 
        n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, 
        n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, 
        n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, 
        n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, 
        n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, 
        n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, 
        n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, 
        n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, 
        n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, 
        n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, 
        n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, 
        n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, 
        n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, 
        n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, 
        n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, 
        n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, 
        n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, 
        n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, 
        n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, 
        n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, 
        n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, 
        n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, 
        n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, 
        n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, 
        n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, 
        n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, 
        n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, 
        n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, 
        n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, 
        n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, 
        n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, 
        n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, 
        n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, 
        n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, 
        n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, 
        n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, 
        n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, 
        n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, 
        n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, 
        n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, 
        n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, 
        n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, 
        n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, 
        n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
        n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, 
        n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, 
        n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, 
        n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, 
        n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, 
        n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, 
        n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, 
        n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, 
        n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, 
        n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, 
        n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, 
        n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, 
        n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, 
        n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, 
        n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, 
        n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, 
        n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, 
        n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, 
        n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, 
        n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, 
        n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, 
        n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, 
        n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, 
        n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, 
        n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, 
        n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, 
        n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, 
        n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, 
        n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, 
        n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, 
        n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, 
        n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, 
        n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, 
        n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, 
        n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, 
        n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, 
        n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, 
        n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, 
        n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, 
        n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, 
        n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, 
        n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, 
        n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, 
        n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, 
        n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, 
        n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, 
        n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, 
        n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, 
        n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, 
        n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, 
        n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, 
        n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, 
        n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, 
        n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, 
        n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, 
        n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, 
        n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, 
        n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, 
        n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, 
        n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, 
        n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, 
        n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, 
        n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, 
        n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, 
        n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, 
        n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, 
        n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, 
        n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, 
        n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, 
        n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, 
        n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, 
        n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, 
        n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, 
        n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, 
        n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, 
        n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, 
        n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, 
        n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, 
        n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, 
        n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, 
        n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, 
        n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, 
        n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, 
        n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, 
        n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, 
        n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, 
        n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, 
        n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, 
        n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, 
        n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, 
        n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, 
        n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, 
        n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, 
        n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, 
        n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, 
        n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, 
        n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, 
        n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, 
        n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, 
        n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, 
        n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, 
        n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, 
        n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, 
        n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, 
        n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, 
        n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, 
        n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, 
        n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, 
        n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, 
        n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, 
        n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, 
        n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, 
        n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, 
        n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, 
        n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, 
        n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, 
        n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, 
        n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, 
        n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, 
        n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, 
        n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, 
        n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, 
        n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, 
        n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, 
        n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, 
        n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, 
        n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, 
        n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, 
        n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, 
        n4255, n4256, n4257, n4258, n4259, n4260, n4262, n4263, 
        n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, 
        n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, 
        n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, 
        n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, 
        n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, 
        n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, 
        n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, 
        n4320, n4321, n4322, n4323, n4324, n4325;
    
    Mux_5u_32u Mux_3 (.sel({ra0}), .data({pcout[31], spout[31], lrout[31], 
            stout[31], \regs[27] [31], \regs[26] [31], \regs[25] [31], 
            \regs[24] [31], \regs[23] [31], \regs[22] [31], \regs[21] [31], 
            \regs[20] [31], \regs[19] [31], \regs[18] [31], \regs[17] [31], 
            \regs[16] [31], \regs[15] [31], \regs[14] [31], \regs[13] [31], 
            \regs[12] [31], \regs[11] [31], \regs[10] [31], \regs[9] [31], 
            \regs[8] [31], \regs[7] [31], \regs[6] [31], \regs[5] [31], 
            \regs[4] [31], \regs[3] [31], \regs[2] [31], \regs[1] [31], 
            \regs[0] [31]}), .o(rd0[31]));   // regs.v(30)
    Mux_5u_32u Mux_4 (.sel({ra0}), .data({pcout[30], spout[30], lrout[30], 
            stout[30], \regs[27] [30], \regs[26] [30], \regs[25] [30], 
            \regs[24] [30], \regs[23] [30], \regs[22] [30], \regs[21] [30], 
            \regs[20] [30], \regs[19] [30], \regs[18] [30], \regs[17] [30], 
            \regs[16] [30], \regs[15] [30], \regs[14] [30], \regs[13] [30], 
            \regs[12] [30], \regs[11] [30], \regs[10] [30], \regs[9] [30], 
            \regs[8] [30], \regs[7] [30], \regs[6] [30], \regs[5] [30], 
            \regs[4] [30], \regs[3] [30], \regs[2] [30], \regs[1] [30], 
            \regs[0] [30]}), .o(rd0[30]));   // regs.v(30)
    Mux_5u_32u Mux_5 (.sel({ra0}), .data({pcout[29], spout[29], lrout[29], 
            stout[29], \regs[27] [29], \regs[26] [29], \regs[25] [29], 
            \regs[24] [29], \regs[23] [29], \regs[22] [29], \regs[21] [29], 
            \regs[20] [29], \regs[19] [29], \regs[18] [29], \regs[17] [29], 
            \regs[16] [29], \regs[15] [29], \regs[14] [29], \regs[13] [29], 
            \regs[12] [29], \regs[11] [29], \regs[10] [29], \regs[9] [29], 
            \regs[8] [29], \regs[7] [29], \regs[6] [29], \regs[5] [29], 
            \regs[4] [29], \regs[3] [29], \regs[2] [29], \regs[1] [29], 
            \regs[0] [29]}), .o(rd0[29]));   // regs.v(30)
    Mux_5u_32u Mux_6 (.sel({ra0}), .data({pcout[28], spout[28], lrout[28], 
            stout[28], \regs[27] [28], \regs[26] [28], \regs[25] [28], 
            \regs[24] [28], \regs[23] [28], \regs[22] [28], \regs[21] [28], 
            \regs[20] [28], \regs[19] [28], \regs[18] [28], \regs[17] [28], 
            \regs[16] [28], \regs[15] [28], \regs[14] [28], \regs[13] [28], 
            \regs[12] [28], \regs[11] [28], \regs[10] [28], \regs[9] [28], 
            \regs[8] [28], \regs[7] [28], \regs[6] [28], \regs[5] [28], 
            \regs[4] [28], \regs[3] [28], \regs[2] [28], \regs[1] [28], 
            \regs[0] [28]}), .o(rd0[28]));   // regs.v(30)
    Mux_5u_32u Mux_7 (.sel({ra0}), .data({pcout[27], spout[27], lrout[27], 
            stout[27], \regs[27] [27], \regs[26] [27], \regs[25] [27], 
            \regs[24] [27], \regs[23] [27], \regs[22] [27], \regs[21] [27], 
            \regs[20] [27], \regs[19] [27], \regs[18] [27], \regs[17] [27], 
            \regs[16] [27], \regs[15] [27], \regs[14] [27], \regs[13] [27], 
            \regs[12] [27], \regs[11] [27], \regs[10] [27], \regs[9] [27], 
            \regs[8] [27], \regs[7] [27], \regs[6] [27], \regs[5] [27], 
            \regs[4] [27], \regs[3] [27], \regs[2] [27], \regs[1] [27], 
            \regs[0] [27]}), .o(rd0[27]));   // regs.v(30)
    Mux_5u_32u Mux_8 (.sel({ra0}), .data({pcout[26], spout[26], lrout[26], 
            stout[26], \regs[27] [26], \regs[26] [26], \regs[25] [26], 
            \regs[24] [26], \regs[23] [26], \regs[22] [26], \regs[21] [26], 
            \regs[20] [26], \regs[19] [26], \regs[18] [26], \regs[17] [26], 
            \regs[16] [26], \regs[15] [26], \regs[14] [26], \regs[13] [26], 
            \regs[12] [26], \regs[11] [26], \regs[10] [26], \regs[9] [26], 
            \regs[8] [26], \regs[7] [26], \regs[6] [26], \regs[5] [26], 
            \regs[4] [26], \regs[3] [26], \regs[2] [26], \regs[1] [26], 
            \regs[0] [26]}), .o(rd0[26]));   // regs.v(30)
    Mux_5u_32u Mux_9 (.sel({ra0}), .data({pcout[25], spout[25], lrout[25], 
            stout[25], \regs[27] [25], \regs[26] [25], \regs[25] [25], 
            \regs[24] [25], \regs[23] [25], \regs[22] [25], \regs[21] [25], 
            \regs[20] [25], \regs[19] [25], \regs[18] [25], \regs[17] [25], 
            \regs[16] [25], \regs[15] [25], \regs[14] [25], \regs[13] [25], 
            \regs[12] [25], \regs[11] [25], \regs[10] [25], \regs[9] [25], 
            \regs[8] [25], \regs[7] [25], \regs[6] [25], \regs[5] [25], 
            \regs[4] [25], \regs[3] [25], \regs[2] [25], \regs[1] [25], 
            \regs[0] [25]}), .o(rd0[25]));   // regs.v(30)
    Mux_5u_32u Mux_10 (.sel({ra0}), .data({pcout[24], spout[24], lrout[24], 
            stout[24], \regs[27] [24], \regs[26] [24], \regs[25] [24], 
            \regs[24] [24], \regs[23] [24], \regs[22] [24], \regs[21] [24], 
            \regs[20] [24], \regs[19] [24], \regs[18] [24], \regs[17] [24], 
            \regs[16] [24], \regs[15] [24], \regs[14] [24], \regs[13] [24], 
            \regs[12] [24], \regs[11] [24], \regs[10] [24], \regs[9] [24], 
            \regs[8] [24], \regs[7] [24], \regs[6] [24], \regs[5] [24], 
            \regs[4] [24], \regs[3] [24], \regs[2] [24], \regs[1] [24], 
            \regs[0] [24]}), .o(rd0[24]));   // regs.v(30)
    Mux_5u_32u Mux_11 (.sel({ra0}), .data({pcout[23], spout[23], lrout[23], 
            stout[23], \regs[27] [23], \regs[26] [23], \regs[25] [23], 
            \regs[24] [23], \regs[23] [23], \regs[22] [23], \regs[21] [23], 
            \regs[20] [23], \regs[19] [23], \regs[18] [23], \regs[17] [23], 
            \regs[16] [23], \regs[15] [23], \regs[14] [23], \regs[13] [23], 
            \regs[12] [23], \regs[11] [23], \regs[10] [23], \regs[9] [23], 
            \regs[8] [23], \regs[7] [23], \regs[6] [23], \regs[5] [23], 
            \regs[4] [23], \regs[3] [23], \regs[2] [23], \regs[1] [23], 
            \regs[0] [23]}), .o(rd0[23]));   // regs.v(30)
    Mux_5u_32u Mux_12 (.sel({ra0}), .data({pcout[22], spout[22], lrout[22], 
            stout[22], \regs[27] [22], \regs[26] [22], \regs[25] [22], 
            \regs[24] [22], \regs[23] [22], \regs[22] [22], \regs[21] [22], 
            \regs[20] [22], \regs[19] [22], \regs[18] [22], \regs[17] [22], 
            \regs[16] [22], \regs[15] [22], \regs[14] [22], \regs[13] [22], 
            \regs[12] [22], \regs[11] [22], \regs[10] [22], \regs[9] [22], 
            \regs[8] [22], \regs[7] [22], \regs[6] [22], \regs[5] [22], 
            \regs[4] [22], \regs[3] [22], \regs[2] [22], \regs[1] [22], 
            \regs[0] [22]}), .o(rd0[22]));   // regs.v(30)
    Mux_5u_32u Mux_13 (.sel({ra0}), .data({pcout[21], spout[21], lrout[21], 
            stout[21], \regs[27] [21], \regs[26] [21], \regs[25] [21], 
            \regs[24] [21], \regs[23] [21], \regs[22] [21], \regs[21] [21], 
            \regs[20] [21], \regs[19] [21], \regs[18] [21], \regs[17] [21], 
            \regs[16] [21], \regs[15] [21], \regs[14] [21], \regs[13] [21], 
            \regs[12] [21], \regs[11] [21], \regs[10] [21], \regs[9] [21], 
            \regs[8] [21], \regs[7] [21], \regs[6] [21], \regs[5] [21], 
            \regs[4] [21], \regs[3] [21], \regs[2] [21], \regs[1] [21], 
            \regs[0] [21]}), .o(rd0[21]));   // regs.v(30)
    Mux_5u_32u Mux_14 (.sel({ra0}), .data({pcout[20], spout[20], lrout[20], 
            stout[20], \regs[27] [20], \regs[26] [20], \regs[25] [20], 
            \regs[24] [20], \regs[23] [20], \regs[22] [20], \regs[21] [20], 
            \regs[20] [20], \regs[19] [20], \regs[18] [20], \regs[17] [20], 
            \regs[16] [20], \regs[15] [20], \regs[14] [20], \regs[13] [20], 
            \regs[12] [20], \regs[11] [20], \regs[10] [20], \regs[9] [20], 
            \regs[8] [20], \regs[7] [20], \regs[6] [20], \regs[5] [20], 
            \regs[4] [20], \regs[3] [20], \regs[2] [20], \regs[1] [20], 
            \regs[0] [20]}), .o(rd0[20]));   // regs.v(30)
    Mux_5u_32u Mux_15 (.sel({ra0}), .data({pcout[19], spout[19], lrout[19], 
            stout[19], \regs[27] [19], \regs[26] [19], \regs[25] [19], 
            \regs[24] [19], \regs[23] [19], \regs[22] [19], \regs[21] [19], 
            \regs[20] [19], \regs[19] [19], \regs[18] [19], \regs[17] [19], 
            \regs[16] [19], \regs[15] [19], \regs[14] [19], \regs[13] [19], 
            \regs[12] [19], \regs[11] [19], \regs[10] [19], \regs[9] [19], 
            \regs[8] [19], \regs[7] [19], \regs[6] [19], \regs[5] [19], 
            \regs[4] [19], \regs[3] [19], \regs[2] [19], \regs[1] [19], 
            \regs[0] [19]}), .o(rd0[19]));   // regs.v(30)
    Mux_5u_32u Mux_16 (.sel({ra0}), .data({pcout[18], spout[18], lrout[18], 
            stout[18], \regs[27] [18], \regs[26] [18], \regs[25] [18], 
            \regs[24] [18], \regs[23] [18], \regs[22] [18], \regs[21] [18], 
            \regs[20] [18], \regs[19] [18], \regs[18] [18], \regs[17] [18], 
            \regs[16] [18], \regs[15] [18], \regs[14] [18], \regs[13] [18], 
            \regs[12] [18], \regs[11] [18], \regs[10] [18], \regs[9] [18], 
            \regs[8] [18], \regs[7] [18], \regs[6] [18], \regs[5] [18], 
            \regs[4] [18], \regs[3] [18], \regs[2] [18], \regs[1] [18], 
            \regs[0] [18]}), .o(rd0[18]));   // regs.v(30)
    Mux_5u_32u Mux_17 (.sel({ra0}), .data({pcout[17], spout[17], lrout[17], 
            stout[17], \regs[27] [17], \regs[26] [17], \regs[25] [17], 
            \regs[24] [17], \regs[23] [17], \regs[22] [17], \regs[21] [17], 
            \regs[20] [17], \regs[19] [17], \regs[18] [17], \regs[17] [17], 
            \regs[16] [17], \regs[15] [17], \regs[14] [17], \regs[13] [17], 
            \regs[12] [17], \regs[11] [17], \regs[10] [17], \regs[9] [17], 
            \regs[8] [17], \regs[7] [17], \regs[6] [17], \regs[5] [17], 
            \regs[4] [17], \regs[3] [17], \regs[2] [17], \regs[1] [17], 
            \regs[0] [17]}), .o(rd0[17]));   // regs.v(30)
    Mux_5u_32u Mux_18 (.sel({ra0}), .data({pcout[16], spout[16], lrout[16], 
            stout[16], \regs[27] [16], \regs[26] [16], \regs[25] [16], 
            \regs[24] [16], \regs[23] [16], \regs[22] [16], \regs[21] [16], 
            \regs[20] [16], \regs[19] [16], \regs[18] [16], \regs[17] [16], 
            \regs[16] [16], \regs[15] [16], \regs[14] [16], \regs[13] [16], 
            \regs[12] [16], \regs[11] [16], \regs[10] [16], \regs[9] [16], 
            \regs[8] [16], \regs[7] [16], \regs[6] [16], \regs[5] [16], 
            \regs[4] [16], \regs[3] [16], \regs[2] [16], \regs[1] [16], 
            \regs[0] [16]}), .o(rd0[16]));   // regs.v(30)
    Mux_5u_32u Mux_19 (.sel({ra0}), .data({pcout[15], spout[15], lrout[15], 
            stout[15], \regs[27] [15], \regs[26] [15], \regs[25] [15], 
            \regs[24] [15], \regs[23] [15], \regs[22] [15], \regs[21] [15], 
            \regs[20] [15], \regs[19] [15], \regs[18] [15], \regs[17] [15], 
            \regs[16] [15], \regs[15] [15], \regs[14] [15], \regs[13] [15], 
            \regs[12] [15], \regs[11] [15], \regs[10] [15], \regs[9] [15], 
            \regs[8] [15], \regs[7] [15], \regs[6] [15], \regs[5] [15], 
            \regs[4] [15], \regs[3] [15], \regs[2] [15], \regs[1] [15], 
            \regs[0] [15]}), .o(rd0[15]));   // regs.v(30)
    Mux_5u_32u Mux_20 (.sel({ra0}), .data({pcout[14], spout[14], lrout[14], 
            stout[14], \regs[27] [14], \regs[26] [14], \regs[25] [14], 
            \regs[24] [14], \regs[23] [14], \regs[22] [14], \regs[21] [14], 
            \regs[20] [14], \regs[19] [14], \regs[18] [14], \regs[17] [14], 
            \regs[16] [14], \regs[15] [14], \regs[14] [14], \regs[13] [14], 
            \regs[12] [14], \regs[11] [14], \regs[10] [14], \regs[9] [14], 
            \regs[8] [14], \regs[7] [14], \regs[6] [14], \regs[5] [14], 
            \regs[4] [14], \regs[3] [14], \regs[2] [14], \regs[1] [14], 
            \regs[0] [14]}), .o(rd0[14]));   // regs.v(30)
    Mux_5u_32u Mux_21 (.sel({ra0}), .data({pcout[13], spout[13], lrout[13], 
            stout[13], \regs[27] [13], \regs[26] [13], \regs[25] [13], 
            \regs[24] [13], \regs[23] [13], \regs[22] [13], \regs[21] [13], 
            \regs[20] [13], \regs[19] [13], \regs[18] [13], \regs[17] [13], 
            \regs[16] [13], \regs[15] [13], \regs[14] [13], \regs[13] [13], 
            \regs[12] [13], \regs[11] [13], \regs[10] [13], \regs[9] [13], 
            \regs[8] [13], \regs[7] [13], \regs[6] [13], \regs[5] [13], 
            \regs[4] [13], \regs[3] [13], \regs[2] [13], \regs[1] [13], 
            \regs[0] [13]}), .o(rd0[13]));   // regs.v(30)
    Mux_5u_32u Mux_22 (.sel({ra0}), .data({pcout[12], spout[12], lrout[12], 
            stout[12], \regs[27] [12], \regs[26] [12], \regs[25] [12], 
            \regs[24] [12], \regs[23] [12], \regs[22] [12], \regs[21] [12], 
            \regs[20] [12], \regs[19] [12], \regs[18] [12], \regs[17] [12], 
            \regs[16] [12], \regs[15] [12], \regs[14] [12], \regs[13] [12], 
            \regs[12] [12], \regs[11] [12], \regs[10] [12], \regs[9] [12], 
            \regs[8] [12], \regs[7] [12], \regs[6] [12], \regs[5] [12], 
            \regs[4] [12], \regs[3] [12], \regs[2] [12], \regs[1] [12], 
            \regs[0] [12]}), .o(rd0[12]));   // regs.v(30)
    Mux_5u_32u Mux_23 (.sel({ra0}), .data({pcout[11], spout[11], lrout[11], 
            stout[11], \regs[27] [11], \regs[26] [11], \regs[25] [11], 
            \regs[24] [11], \regs[23] [11], \regs[22] [11], \regs[21] [11], 
            \regs[20] [11], \regs[19] [11], \regs[18] [11], \regs[17] [11], 
            \regs[16] [11], \regs[15] [11], \regs[14] [11], \regs[13] [11], 
            \regs[12] [11], \regs[11] [11], \regs[10] [11], \regs[9] [11], 
            \regs[8] [11], \regs[7] [11], \regs[6] [11], \regs[5] [11], 
            \regs[4] [11], \regs[3] [11], \regs[2] [11], \regs[1] [11], 
            \regs[0] [11]}), .o(rd0[11]));   // regs.v(30)
    Mux_5u_32u Mux_24 (.sel({ra0}), .data({pcout[10], spout[10], lrout[10], 
            stout[10], \regs[27] [10], \regs[26] [10], \regs[25] [10], 
            \regs[24] [10], \regs[23] [10], \regs[22] [10], \regs[21] [10], 
            \regs[20] [10], \regs[19] [10], \regs[18] [10], \regs[17] [10], 
            \regs[16] [10], \regs[15] [10], \regs[14] [10], \regs[13] [10], 
            \regs[12] [10], \regs[11] [10], \regs[10] [10], \regs[9] [10], 
            \regs[8] [10], \regs[7] [10], \regs[6] [10], \regs[5] [10], 
            \regs[4] [10], \regs[3] [10], \regs[2] [10], \regs[1] [10], 
            \regs[0] [10]}), .o(rd0[10]));   // regs.v(30)
    Mux_5u_32u Mux_25 (.sel({ra0}), .data({pcout[9], spout[9], lrout[9], 
            stout[9], \regs[27] [9], \regs[26] [9], \regs[25] [9], \regs[24] [9], 
            \regs[23] [9], \regs[22] [9], \regs[21] [9], \regs[20] [9], 
            \regs[19] [9], \regs[18] [9], \regs[17] [9], \regs[16] [9], 
            \regs[15] [9], \regs[14] [9], \regs[13] [9], \regs[12] [9], 
            \regs[11] [9], \regs[10] [9], \regs[9] [9], \regs[8] [9], 
            \regs[7] [9], \regs[6] [9], \regs[5] [9], \regs[4] [9], 
            \regs[3] [9], \regs[2] [9], \regs[1] [9], \regs[0] [9]}), 
            .o(rd0[9]));   // regs.v(30)
    Mux_5u_32u Mux_26 (.sel({ra0}), .data({pcout[8], spout[8], lrout[8], 
            stout[8], \regs[27] [8], \regs[26] [8], \regs[25] [8], \regs[24] [8], 
            \regs[23] [8], \regs[22] [8], \regs[21] [8], \regs[20] [8], 
            \regs[19] [8], \regs[18] [8], \regs[17] [8], \regs[16] [8], 
            \regs[15] [8], \regs[14] [8], \regs[13] [8], \regs[12] [8], 
            \regs[11] [8], \regs[10] [8], \regs[9] [8], \regs[8] [8], 
            \regs[7] [8], \regs[6] [8], \regs[5] [8], \regs[4] [8], 
            \regs[3] [8], \regs[2] [8], \regs[1] [8], \regs[0] [8]}), 
            .o(rd0[8]));   // regs.v(30)
    Mux_5u_32u Mux_27 (.sel({ra0}), .data({pcout[7], spout[7], lrout[7], 
            stout[7], \regs[27] [7], \regs[26] [7], \regs[25] [7], \regs[24] [7], 
            \regs[23] [7], \regs[22] [7], \regs[21] [7], \regs[20] [7], 
            \regs[19] [7], \regs[18] [7], \regs[17] [7], \regs[16] [7], 
            \regs[15] [7], \regs[14] [7], \regs[13] [7], \regs[12] [7], 
            \regs[11] [7], \regs[10] [7], \regs[9] [7], \regs[8] [7], 
            \regs[7] [7], \regs[6] [7], \regs[5] [7], \regs[4] [7], 
            \regs[3] [7], \regs[2] [7], \regs[1] [7], \regs[0] [7]}), 
            .o(rd0[7]));   // regs.v(30)
    Mux_5u_32u Mux_28 (.sel({ra0}), .data({pcout[6], spout[6], lrout[6], 
            stout[6], \regs[27] [6], \regs[26] [6], \regs[25] [6], \regs[24] [6], 
            \regs[23] [6], \regs[22] [6], \regs[21] [6], \regs[20] [6], 
            \regs[19] [6], \regs[18] [6], \regs[17] [6], \regs[16] [6], 
            \regs[15] [6], \regs[14] [6], \regs[13] [6], \regs[12] [6], 
            \regs[11] [6], \regs[10] [6], \regs[9] [6], \regs[8] [6], 
            \regs[7] [6], \regs[6] [6], \regs[5] [6], \regs[4] [6], 
            \regs[3] [6], \regs[2] [6], \regs[1] [6], \regs[0] [6]}), 
            .o(rd0[6]));   // regs.v(30)
    Mux_5u_32u Mux_29 (.sel({ra0}), .data({pcout[5], spout[5], lrout[5], 
            stout[5], \regs[27] [5], \regs[26] [5], \regs[25] [5], \regs[24] [5], 
            \regs[23] [5], \regs[22] [5], \regs[21] [5], \regs[20] [5], 
            \regs[19] [5], \regs[18] [5], \regs[17] [5], \regs[16] [5], 
            \regs[15] [5], \regs[14] [5], \regs[13] [5], \regs[12] [5], 
            \regs[11] [5], \regs[10] [5], \regs[9] [5], \regs[8] [5], 
            \regs[7] [5], \regs[6] [5], \regs[5] [5], \regs[4] [5], 
            \regs[3] [5], \regs[2] [5], \regs[1] [5], \regs[0] [5]}), 
            .o(rd0[5]));   // regs.v(30)
    Mux_5u_32u Mux_30 (.sel({ra0}), .data({pcout[4], spout[4], lrout[4], 
            stout[4], \regs[27] [4], \regs[26] [4], \regs[25] [4], \regs[24] [4], 
            \regs[23] [4], \regs[22] [4], \regs[21] [4], \regs[20] [4], 
            \regs[19] [4], \regs[18] [4], \regs[17] [4], \regs[16] [4], 
            \regs[15] [4], \regs[14] [4], \regs[13] [4], \regs[12] [4], 
            \regs[11] [4], \regs[10] [4], \regs[9] [4], \regs[8] [4], 
            \regs[7] [4], \regs[6] [4], \regs[5] [4], \regs[4] [4], 
            \regs[3] [4], \regs[2] [4], \regs[1] [4], \regs[0] [4]}), 
            .o(rd0[4]));   // regs.v(30)
    Mux_5u_32u Mux_31 (.sel({ra0}), .data({pcout[3], spout[3], lrout[3], 
            stout[3], \regs[27] [3], \regs[26] [3], \regs[25] [3], \regs[24] [3], 
            \regs[23] [3], \regs[22] [3], \regs[21] [3], \regs[20] [3], 
            \regs[19] [3], \regs[18] [3], \regs[17] [3], \regs[16] [3], 
            \regs[15] [3], \regs[14] [3], \regs[13] [3], \regs[12] [3], 
            \regs[11] [3], \regs[10] [3], \regs[9] [3], \regs[8] [3], 
            \regs[7] [3], \regs[6] [3], \regs[5] [3], \regs[4] [3], 
            \regs[3] [3], \regs[2] [3], \regs[1] [3], \regs[0] [3]}), 
            .o(rd0[3]));   // regs.v(30)
    Mux_5u_32u Mux_32 (.sel({ra0}), .data({pcout[2], spout[2], lrout[2], 
            stout[2], \regs[27] [2], \regs[26] [2], \regs[25] [2], \regs[24] [2], 
            \regs[23] [2], \regs[22] [2], \regs[21] [2], \regs[20] [2], 
            \regs[19] [2], \regs[18] [2], \regs[17] [2], \regs[16] [2], 
            \regs[15] [2], \regs[14] [2], \regs[13] [2], \regs[12] [2], 
            \regs[11] [2], \regs[10] [2], \regs[9] [2], \regs[8] [2], 
            \regs[7] [2], \regs[6] [2], \regs[5] [2], \regs[4] [2], 
            \regs[3] [2], \regs[2] [2], \regs[1] [2], \regs[0] [2]}), 
            .o(rd0[2]));   // regs.v(30)
    Mux_5u_32u Mux_33 (.sel({ra0}), .data({pcout[1], spout[1], lrout[1], 
            stout[1], \regs[27] [1], \regs[26] [1], \regs[25] [1], \regs[24] [1], 
            \regs[23] [1], \regs[22] [1], \regs[21] [1], \regs[20] [1], 
            \regs[19] [1], \regs[18] [1], \regs[17] [1], \regs[16] [1], 
            \regs[15] [1], \regs[14] [1], \regs[13] [1], \regs[12] [1], 
            \regs[11] [1], \regs[10] [1], \regs[9] [1], \regs[8] [1], 
            \regs[7] [1], \regs[6] [1], \regs[5] [1], \regs[4] [1], 
            \regs[3] [1], \regs[2] [1], \regs[1] [1], \regs[0] [1]}), 
            .o(rd0[1]));   // regs.v(30)
    Mux_5u_32u Mux_34 (.sel({ra0}), .data({pcout[0], spout[0], lrout[0], 
            stout[0], \regs[27] [0], \regs[26] [0], \regs[25] [0], \regs[24] [0], 
            \regs[23] [0], \regs[22] [0], \regs[21] [0], \regs[20] [0], 
            \regs[19] [0], \regs[18] [0], \regs[17] [0], \regs[16] [0], 
            \regs[15] [0], \regs[14] [0], \regs[13] [0], \regs[12] [0], 
            \regs[11] [0], \regs[10] [0], \regs[9] [0], \regs[8] [0], 
            \regs[7] [0], \regs[6] [0], \regs[5] [0], \regs[4] [0], 
            \regs[3] [0], \regs[2] [0], \regs[1] [0], \regs[0] [0]}), 
            .o(rd0[0]));   // regs.v(30)
    Mux_5u_32u Mux_35 (.sel({ra1}), .data({pcout[31], spout[31], lrout[31], 
            stout[31], \regs[27] [31], \regs[26] [31], \regs[25] [31], 
            \regs[24] [31], \regs[23] [31], \regs[22] [31], \regs[21] [31], 
            \regs[20] [31], \regs[19] [31], \regs[18] [31], \regs[17] [31], 
            \regs[16] [31], \regs[15] [31], \regs[14] [31], \regs[13] [31], 
            \regs[12] [31], \regs[11] [31], \regs[10] [31], \regs[9] [31], 
            \regs[8] [31], \regs[7] [31], \regs[6] [31], \regs[5] [31], 
            \regs[4] [31], \regs[3] [31], \regs[2] [31], \regs[1] [31], 
            \regs[0] [31]}), .o(rd1[31]));   // regs.v(31)
    Mux_5u_32u Mux_36 (.sel({ra1}), .data({pcout[30], spout[30], lrout[30], 
            stout[30], \regs[27] [30], \regs[26] [30], \regs[25] [30], 
            \regs[24] [30], \regs[23] [30], \regs[22] [30], \regs[21] [30], 
            \regs[20] [30], \regs[19] [30], \regs[18] [30], \regs[17] [30], 
            \regs[16] [30], \regs[15] [30], \regs[14] [30], \regs[13] [30], 
            \regs[12] [30], \regs[11] [30], \regs[10] [30], \regs[9] [30], 
            \regs[8] [30], \regs[7] [30], \regs[6] [30], \regs[5] [30], 
            \regs[4] [30], \regs[3] [30], \regs[2] [30], \regs[1] [30], 
            \regs[0] [30]}), .o(rd1[30]));   // regs.v(31)
    Mux_5u_32u Mux_37 (.sel({ra1}), .data({pcout[29], spout[29], lrout[29], 
            stout[29], \regs[27] [29], \regs[26] [29], \regs[25] [29], 
            \regs[24] [29], \regs[23] [29], \regs[22] [29], \regs[21] [29], 
            \regs[20] [29], \regs[19] [29], \regs[18] [29], \regs[17] [29], 
            \regs[16] [29], \regs[15] [29], \regs[14] [29], \regs[13] [29], 
            \regs[12] [29], \regs[11] [29], \regs[10] [29], \regs[9] [29], 
            \regs[8] [29], \regs[7] [29], \regs[6] [29], \regs[5] [29], 
            \regs[4] [29], \regs[3] [29], \regs[2] [29], \regs[1] [29], 
            \regs[0] [29]}), .o(rd1[29]));   // regs.v(31)
    Mux_5u_32u Mux_38 (.sel({ra1}), .data({pcout[28], spout[28], lrout[28], 
            stout[28], \regs[27] [28], \regs[26] [28], \regs[25] [28], 
            \regs[24] [28], \regs[23] [28], \regs[22] [28], \regs[21] [28], 
            \regs[20] [28], \regs[19] [28], \regs[18] [28], \regs[17] [28], 
            \regs[16] [28], \regs[15] [28], \regs[14] [28], \regs[13] [28], 
            \regs[12] [28], \regs[11] [28], \regs[10] [28], \regs[9] [28], 
            \regs[8] [28], \regs[7] [28], \regs[6] [28], \regs[5] [28], 
            \regs[4] [28], \regs[3] [28], \regs[2] [28], \regs[1] [28], 
            \regs[0] [28]}), .o(rd1[28]));   // regs.v(31)
    Mux_5u_32u Mux_39 (.sel({ra1}), .data({pcout[27], spout[27], lrout[27], 
            stout[27], \regs[27] [27], \regs[26] [27], \regs[25] [27], 
            \regs[24] [27], \regs[23] [27], \regs[22] [27], \regs[21] [27], 
            \regs[20] [27], \regs[19] [27], \regs[18] [27], \regs[17] [27], 
            \regs[16] [27], \regs[15] [27], \regs[14] [27], \regs[13] [27], 
            \regs[12] [27], \regs[11] [27], \regs[10] [27], \regs[9] [27], 
            \regs[8] [27], \regs[7] [27], \regs[6] [27], \regs[5] [27], 
            \regs[4] [27], \regs[3] [27], \regs[2] [27], \regs[1] [27], 
            \regs[0] [27]}), .o(rd1[27]));   // regs.v(31)
    Mux_5u_32u Mux_40 (.sel({ra1}), .data({pcout[26], spout[26], lrout[26], 
            stout[26], \regs[27] [26], \regs[26] [26], \regs[25] [26], 
            \regs[24] [26], \regs[23] [26], \regs[22] [26], \regs[21] [26], 
            \regs[20] [26], \regs[19] [26], \regs[18] [26], \regs[17] [26], 
            \regs[16] [26], \regs[15] [26], \regs[14] [26], \regs[13] [26], 
            \regs[12] [26], \regs[11] [26], \regs[10] [26], \regs[9] [26], 
            \regs[8] [26], \regs[7] [26], \regs[6] [26], \regs[5] [26], 
            \regs[4] [26], \regs[3] [26], \regs[2] [26], \regs[1] [26], 
            \regs[0] [26]}), .o(rd1[26]));   // regs.v(31)
    Mux_5u_32u Mux_41 (.sel({ra1}), .data({pcout[25], spout[25], lrout[25], 
            stout[25], \regs[27] [25], \regs[26] [25], \regs[25] [25], 
            \regs[24] [25], \regs[23] [25], \regs[22] [25], \regs[21] [25], 
            \regs[20] [25], \regs[19] [25], \regs[18] [25], \regs[17] [25], 
            \regs[16] [25], \regs[15] [25], \regs[14] [25], \regs[13] [25], 
            \regs[12] [25], \regs[11] [25], \regs[10] [25], \regs[9] [25], 
            \regs[8] [25], \regs[7] [25], \regs[6] [25], \regs[5] [25], 
            \regs[4] [25], \regs[3] [25], \regs[2] [25], \regs[1] [25], 
            \regs[0] [25]}), .o(rd1[25]));   // regs.v(31)
    Mux_5u_32u Mux_42 (.sel({ra1}), .data({pcout[24], spout[24], lrout[24], 
            stout[24], \regs[27] [24], \regs[26] [24], \regs[25] [24], 
            \regs[24] [24], \regs[23] [24], \regs[22] [24], \regs[21] [24], 
            \regs[20] [24], \regs[19] [24], \regs[18] [24], \regs[17] [24], 
            \regs[16] [24], \regs[15] [24], \regs[14] [24], \regs[13] [24], 
            \regs[12] [24], \regs[11] [24], \regs[10] [24], \regs[9] [24], 
            \regs[8] [24], \regs[7] [24], \regs[6] [24], \regs[5] [24], 
            \regs[4] [24], \regs[3] [24], \regs[2] [24], \regs[1] [24], 
            \regs[0] [24]}), .o(rd1[24]));   // regs.v(31)
    Mux_5u_32u Mux_43 (.sel({ra1}), .data({pcout[23], spout[23], lrout[23], 
            stout[23], \regs[27] [23], \regs[26] [23], \regs[25] [23], 
            \regs[24] [23], \regs[23] [23], \regs[22] [23], \regs[21] [23], 
            \regs[20] [23], \regs[19] [23], \regs[18] [23], \regs[17] [23], 
            \regs[16] [23], \regs[15] [23], \regs[14] [23], \regs[13] [23], 
            \regs[12] [23], \regs[11] [23], \regs[10] [23], \regs[9] [23], 
            \regs[8] [23], \regs[7] [23], \regs[6] [23], \regs[5] [23], 
            \regs[4] [23], \regs[3] [23], \regs[2] [23], \regs[1] [23], 
            \regs[0] [23]}), .o(rd1[23]));   // regs.v(31)
    Mux_5u_32u Mux_44 (.sel({ra1}), .data({pcout[22], spout[22], lrout[22], 
            stout[22], \regs[27] [22], \regs[26] [22], \regs[25] [22], 
            \regs[24] [22], \regs[23] [22], \regs[22] [22], \regs[21] [22], 
            \regs[20] [22], \regs[19] [22], \regs[18] [22], \regs[17] [22], 
            \regs[16] [22], \regs[15] [22], \regs[14] [22], \regs[13] [22], 
            \regs[12] [22], \regs[11] [22], \regs[10] [22], \regs[9] [22], 
            \regs[8] [22], \regs[7] [22], \regs[6] [22], \regs[5] [22], 
            \regs[4] [22], \regs[3] [22], \regs[2] [22], \regs[1] [22], 
            \regs[0] [22]}), .o(rd1[22]));   // regs.v(31)
    Mux_5u_32u Mux_45 (.sel({ra1}), .data({pcout[21], spout[21], lrout[21], 
            stout[21], \regs[27] [21], \regs[26] [21], \regs[25] [21], 
            \regs[24] [21], \regs[23] [21], \regs[22] [21], \regs[21] [21], 
            \regs[20] [21], \regs[19] [21], \regs[18] [21], \regs[17] [21], 
            \regs[16] [21], \regs[15] [21], \regs[14] [21], \regs[13] [21], 
            \regs[12] [21], \regs[11] [21], \regs[10] [21], \regs[9] [21], 
            \regs[8] [21], \regs[7] [21], \regs[6] [21], \regs[5] [21], 
            \regs[4] [21], \regs[3] [21], \regs[2] [21], \regs[1] [21], 
            \regs[0] [21]}), .o(rd1[21]));   // regs.v(31)
    Mux_5u_32u Mux_46 (.sel({ra1}), .data({pcout[20], spout[20], lrout[20], 
            stout[20], \regs[27] [20], \regs[26] [20], \regs[25] [20], 
            \regs[24] [20], \regs[23] [20], \regs[22] [20], \regs[21] [20], 
            \regs[20] [20], \regs[19] [20], \regs[18] [20], \regs[17] [20], 
            \regs[16] [20], \regs[15] [20], \regs[14] [20], \regs[13] [20], 
            \regs[12] [20], \regs[11] [20], \regs[10] [20], \regs[9] [20], 
            \regs[8] [20], \regs[7] [20], \regs[6] [20], \regs[5] [20], 
            \regs[4] [20], \regs[3] [20], \regs[2] [20], \regs[1] [20], 
            \regs[0] [20]}), .o(rd1[20]));   // regs.v(31)
    Mux_5u_32u Mux_47 (.sel({ra1}), .data({pcout[19], spout[19], lrout[19], 
            stout[19], \regs[27] [19], \regs[26] [19], \regs[25] [19], 
            \regs[24] [19], \regs[23] [19], \regs[22] [19], \regs[21] [19], 
            \regs[20] [19], \regs[19] [19], \regs[18] [19], \regs[17] [19], 
            \regs[16] [19], \regs[15] [19], \regs[14] [19], \regs[13] [19], 
            \regs[12] [19], \regs[11] [19], \regs[10] [19], \regs[9] [19], 
            \regs[8] [19], \regs[7] [19], \regs[6] [19], \regs[5] [19], 
            \regs[4] [19], \regs[3] [19], \regs[2] [19], \regs[1] [19], 
            \regs[0] [19]}), .o(rd1[19]));   // regs.v(31)
    Mux_5u_32u Mux_48 (.sel({ra1}), .data({pcout[18], spout[18], lrout[18], 
            stout[18], \regs[27] [18], \regs[26] [18], \regs[25] [18], 
            \regs[24] [18], \regs[23] [18], \regs[22] [18], \regs[21] [18], 
            \regs[20] [18], \regs[19] [18], \regs[18] [18], \regs[17] [18], 
            \regs[16] [18], \regs[15] [18], \regs[14] [18], \regs[13] [18], 
            \regs[12] [18], \regs[11] [18], \regs[10] [18], \regs[9] [18], 
            \regs[8] [18], \regs[7] [18], \regs[6] [18], \regs[5] [18], 
            \regs[4] [18], \regs[3] [18], \regs[2] [18], \regs[1] [18], 
            \regs[0] [18]}), .o(rd1[18]));   // regs.v(31)
    Mux_5u_32u Mux_49 (.sel({ra1}), .data({pcout[17], spout[17], lrout[17], 
            stout[17], \regs[27] [17], \regs[26] [17], \regs[25] [17], 
            \regs[24] [17], \regs[23] [17], \regs[22] [17], \regs[21] [17], 
            \regs[20] [17], \regs[19] [17], \regs[18] [17], \regs[17] [17], 
            \regs[16] [17], \regs[15] [17], \regs[14] [17], \regs[13] [17], 
            \regs[12] [17], \regs[11] [17], \regs[10] [17], \regs[9] [17], 
            \regs[8] [17], \regs[7] [17], \regs[6] [17], \regs[5] [17], 
            \regs[4] [17], \regs[3] [17], \regs[2] [17], \regs[1] [17], 
            \regs[0] [17]}), .o(rd1[17]));   // regs.v(31)
    Mux_5u_32u Mux_50 (.sel({ra1}), .data({pcout[16], spout[16], lrout[16], 
            stout[16], \regs[27] [16], \regs[26] [16], \regs[25] [16], 
            \regs[24] [16], \regs[23] [16], \regs[22] [16], \regs[21] [16], 
            \regs[20] [16], \regs[19] [16], \regs[18] [16], \regs[17] [16], 
            \regs[16] [16], \regs[15] [16], \regs[14] [16], \regs[13] [16], 
            \regs[12] [16], \regs[11] [16], \regs[10] [16], \regs[9] [16], 
            \regs[8] [16], \regs[7] [16], \regs[6] [16], \regs[5] [16], 
            \regs[4] [16], \regs[3] [16], \regs[2] [16], \regs[1] [16], 
            \regs[0] [16]}), .o(rd1[16]));   // regs.v(31)
    Mux_5u_32u Mux_51 (.sel({ra1}), .data({pcout[15], spout[15], lrout[15], 
            stout[15], \regs[27] [15], \regs[26] [15], \regs[25] [15], 
            \regs[24] [15], \regs[23] [15], \regs[22] [15], \regs[21] [15], 
            \regs[20] [15], \regs[19] [15], \regs[18] [15], \regs[17] [15], 
            \regs[16] [15], \regs[15] [15], \regs[14] [15], \regs[13] [15], 
            \regs[12] [15], \regs[11] [15], \regs[10] [15], \regs[9] [15], 
            \regs[8] [15], \regs[7] [15], \regs[6] [15], \regs[5] [15], 
            \regs[4] [15], \regs[3] [15], \regs[2] [15], \regs[1] [15], 
            \regs[0] [15]}), .o(rd1[15]));   // regs.v(31)
    Mux_5u_32u Mux_52 (.sel({ra1}), .data({pcout[14], spout[14], lrout[14], 
            stout[14], \regs[27] [14], \regs[26] [14], \regs[25] [14], 
            \regs[24] [14], \regs[23] [14], \regs[22] [14], \regs[21] [14], 
            \regs[20] [14], \regs[19] [14], \regs[18] [14], \regs[17] [14], 
            \regs[16] [14], \regs[15] [14], \regs[14] [14], \regs[13] [14], 
            \regs[12] [14], \regs[11] [14], \regs[10] [14], \regs[9] [14], 
            \regs[8] [14], \regs[7] [14], \regs[6] [14], \regs[5] [14], 
            \regs[4] [14], \regs[3] [14], \regs[2] [14], \regs[1] [14], 
            \regs[0] [14]}), .o(rd1[14]));   // regs.v(31)
    Mux_5u_32u Mux_53 (.sel({ra1}), .data({pcout[13], spout[13], lrout[13], 
            stout[13], \regs[27] [13], \regs[26] [13], \regs[25] [13], 
            \regs[24] [13], \regs[23] [13], \regs[22] [13], \regs[21] [13], 
            \regs[20] [13], \regs[19] [13], \regs[18] [13], \regs[17] [13], 
            \regs[16] [13], \regs[15] [13], \regs[14] [13], \regs[13] [13], 
            \regs[12] [13], \regs[11] [13], \regs[10] [13], \regs[9] [13], 
            \regs[8] [13], \regs[7] [13], \regs[6] [13], \regs[5] [13], 
            \regs[4] [13], \regs[3] [13], \regs[2] [13], \regs[1] [13], 
            \regs[0] [13]}), .o(rd1[13]));   // regs.v(31)
    Mux_5u_32u Mux_54 (.sel({ra1}), .data({pcout[12], spout[12], lrout[12], 
            stout[12], \regs[27] [12], \regs[26] [12], \regs[25] [12], 
            \regs[24] [12], \regs[23] [12], \regs[22] [12], \regs[21] [12], 
            \regs[20] [12], \regs[19] [12], \regs[18] [12], \regs[17] [12], 
            \regs[16] [12], \regs[15] [12], \regs[14] [12], \regs[13] [12], 
            \regs[12] [12], \regs[11] [12], \regs[10] [12], \regs[9] [12], 
            \regs[8] [12], \regs[7] [12], \regs[6] [12], \regs[5] [12], 
            \regs[4] [12], \regs[3] [12], \regs[2] [12], \regs[1] [12], 
            \regs[0] [12]}), .o(rd1[12]));   // regs.v(31)
    Mux_5u_32u Mux_55 (.sel({ra1}), .data({pcout[11], spout[11], lrout[11], 
            stout[11], \regs[27] [11], \regs[26] [11], \regs[25] [11], 
            \regs[24] [11], \regs[23] [11], \regs[22] [11], \regs[21] [11], 
            \regs[20] [11], \regs[19] [11], \regs[18] [11], \regs[17] [11], 
            \regs[16] [11], \regs[15] [11], \regs[14] [11], \regs[13] [11], 
            \regs[12] [11], \regs[11] [11], \regs[10] [11], \regs[9] [11], 
            \regs[8] [11], \regs[7] [11], \regs[6] [11], \regs[5] [11], 
            \regs[4] [11], \regs[3] [11], \regs[2] [11], \regs[1] [11], 
            \regs[0] [11]}), .o(rd1[11]));   // regs.v(31)
    Mux_5u_32u Mux_56 (.sel({ra1}), .data({pcout[10], spout[10], lrout[10], 
            stout[10], \regs[27] [10], \regs[26] [10], \regs[25] [10], 
            \regs[24] [10], \regs[23] [10], \regs[22] [10], \regs[21] [10], 
            \regs[20] [10], \regs[19] [10], \regs[18] [10], \regs[17] [10], 
            \regs[16] [10], \regs[15] [10], \regs[14] [10], \regs[13] [10], 
            \regs[12] [10], \regs[11] [10], \regs[10] [10], \regs[9] [10], 
            \regs[8] [10], \regs[7] [10], \regs[6] [10], \regs[5] [10], 
            \regs[4] [10], \regs[3] [10], \regs[2] [10], \regs[1] [10], 
            \regs[0] [10]}), .o(rd1[10]));   // regs.v(31)
    Mux_5u_32u Mux_57 (.sel({ra1}), .data({pcout[9], spout[9], lrout[9], 
            stout[9], \regs[27] [9], \regs[26] [9], \regs[25] [9], \regs[24] [9], 
            \regs[23] [9], \regs[22] [9], \regs[21] [9], \regs[20] [9], 
            \regs[19] [9], \regs[18] [9], \regs[17] [9], \regs[16] [9], 
            \regs[15] [9], \regs[14] [9], \regs[13] [9], \regs[12] [9], 
            \regs[11] [9], \regs[10] [9], \regs[9] [9], \regs[8] [9], 
            \regs[7] [9], \regs[6] [9], \regs[5] [9], \regs[4] [9], 
            \regs[3] [9], \regs[2] [9], \regs[1] [9], \regs[0] [9]}), 
            .o(rd1[9]));   // regs.v(31)
    Mux_5u_32u Mux_58 (.sel({ra1}), .data({pcout[8], spout[8], lrout[8], 
            stout[8], \regs[27] [8], \regs[26] [8], \regs[25] [8], \regs[24] [8], 
            \regs[23] [8], \regs[22] [8], \regs[21] [8], \regs[20] [8], 
            \regs[19] [8], \regs[18] [8], \regs[17] [8], \regs[16] [8], 
            \regs[15] [8], \regs[14] [8], \regs[13] [8], \regs[12] [8], 
            \regs[11] [8], \regs[10] [8], \regs[9] [8], \regs[8] [8], 
            \regs[7] [8], \regs[6] [8], \regs[5] [8], \regs[4] [8], 
            \regs[3] [8], \regs[2] [8], \regs[1] [8], \regs[0] [8]}), 
            .o(rd1[8]));   // regs.v(31)
    Mux_5u_32u Mux_59 (.sel({ra1}), .data({pcout[7], spout[7], lrout[7], 
            stout[7], \regs[27] [7], \regs[26] [7], \regs[25] [7], \regs[24] [7], 
            \regs[23] [7], \regs[22] [7], \regs[21] [7], \regs[20] [7], 
            \regs[19] [7], \regs[18] [7], \regs[17] [7], \regs[16] [7], 
            \regs[15] [7], \regs[14] [7], \regs[13] [7], \regs[12] [7], 
            \regs[11] [7], \regs[10] [7], \regs[9] [7], \regs[8] [7], 
            \regs[7] [7], \regs[6] [7], \regs[5] [7], \regs[4] [7], 
            \regs[3] [7], \regs[2] [7], \regs[1] [7], \regs[0] [7]}), 
            .o(rd1[7]));   // regs.v(31)
    Mux_5u_32u Mux_60 (.sel({ra1}), .data({pcout[6], spout[6], lrout[6], 
            stout[6], \regs[27] [6], \regs[26] [6], \regs[25] [6], \regs[24] [6], 
            \regs[23] [6], \regs[22] [6], \regs[21] [6], \regs[20] [6], 
            \regs[19] [6], \regs[18] [6], \regs[17] [6], \regs[16] [6], 
            \regs[15] [6], \regs[14] [6], \regs[13] [6], \regs[12] [6], 
            \regs[11] [6], \regs[10] [6], \regs[9] [6], \regs[8] [6], 
            \regs[7] [6], \regs[6] [6], \regs[5] [6], \regs[4] [6], 
            \regs[3] [6], \regs[2] [6], \regs[1] [6], \regs[0] [6]}), 
            .o(rd1[6]));   // regs.v(31)
    Mux_5u_32u Mux_61 (.sel({ra1}), .data({pcout[5], spout[5], lrout[5], 
            stout[5], \regs[27] [5], \regs[26] [5], \regs[25] [5], \regs[24] [5], 
            \regs[23] [5], \regs[22] [5], \regs[21] [5], \regs[20] [5], 
            \regs[19] [5], \regs[18] [5], \regs[17] [5], \regs[16] [5], 
            \regs[15] [5], \regs[14] [5], \regs[13] [5], \regs[12] [5], 
            \regs[11] [5], \regs[10] [5], \regs[9] [5], \regs[8] [5], 
            \regs[7] [5], \regs[6] [5], \regs[5] [5], \regs[4] [5], 
            \regs[3] [5], \regs[2] [5], \regs[1] [5], \regs[0] [5]}), 
            .o(rd1[5]));   // regs.v(31)
    Mux_5u_32u Mux_62 (.sel({ra1}), .data({pcout[4], spout[4], lrout[4], 
            stout[4], \regs[27] [4], \regs[26] [4], \regs[25] [4], \regs[24] [4], 
            \regs[23] [4], \regs[22] [4], \regs[21] [4], \regs[20] [4], 
            \regs[19] [4], \regs[18] [4], \regs[17] [4], \regs[16] [4], 
            \regs[15] [4], \regs[14] [4], \regs[13] [4], \regs[12] [4], 
            \regs[11] [4], \regs[10] [4], \regs[9] [4], \regs[8] [4], 
            \regs[7] [4], \regs[6] [4], \regs[5] [4], \regs[4] [4], 
            \regs[3] [4], \regs[2] [4], \regs[1] [4], \regs[0] [4]}), 
            .o(rd1[4]));   // regs.v(31)
    Mux_5u_32u Mux_63 (.sel({ra1}), .data({pcout[3], spout[3], lrout[3], 
            stout[3], \regs[27] [3], \regs[26] [3], \regs[25] [3], \regs[24] [3], 
            \regs[23] [3], \regs[22] [3], \regs[21] [3], \regs[20] [3], 
            \regs[19] [3], \regs[18] [3], \regs[17] [3], \regs[16] [3], 
            \regs[15] [3], \regs[14] [3], \regs[13] [3], \regs[12] [3], 
            \regs[11] [3], \regs[10] [3], \regs[9] [3], \regs[8] [3], 
            \regs[7] [3], \regs[6] [3], \regs[5] [3], \regs[4] [3], 
            \regs[3] [3], \regs[2] [3], \regs[1] [3], \regs[0] [3]}), 
            .o(rd1[3]));   // regs.v(31)
    Mux_5u_32u Mux_64 (.sel({ra1}), .data({pcout[2], spout[2], lrout[2], 
            stout[2], \regs[27] [2], \regs[26] [2], \regs[25] [2], \regs[24] [2], 
            \regs[23] [2], \regs[22] [2], \regs[21] [2], \regs[20] [2], 
            \regs[19] [2], \regs[18] [2], \regs[17] [2], \regs[16] [2], 
            \regs[15] [2], \regs[14] [2], \regs[13] [2], \regs[12] [2], 
            \regs[11] [2], \regs[10] [2], \regs[9] [2], \regs[8] [2], 
            \regs[7] [2], \regs[6] [2], \regs[5] [2], \regs[4] [2], 
            \regs[3] [2], \regs[2] [2], \regs[1] [2], \regs[0] [2]}), 
            .o(rd1[2]));   // regs.v(31)
    Mux_5u_32u Mux_65 (.sel({ra1}), .data({pcout[1], spout[1], lrout[1], 
            stout[1], \regs[27] [1], \regs[26] [1], \regs[25] [1], \regs[24] [1], 
            \regs[23] [1], \regs[22] [1], \regs[21] [1], \regs[20] [1], 
            \regs[19] [1], \regs[18] [1], \regs[17] [1], \regs[16] [1], 
            \regs[15] [1], \regs[14] [1], \regs[13] [1], \regs[12] [1], 
            \regs[11] [1], \regs[10] [1], \regs[9] [1], \regs[8] [1], 
            \regs[7] [1], \regs[6] [1], \regs[5] [1], \regs[4] [1], 
            \regs[3] [1], \regs[2] [1], \regs[1] [1], \regs[0] [1]}), 
            .o(rd1[1]));   // regs.v(31)
    Mux_5u_32u Mux_66 (.sel({ra1}), .data({pcout[0], spout[0], lrout[0], 
            stout[0], \regs[27] [0], \regs[26] [0], \regs[25] [0], \regs[24] [0], 
            \regs[23] [0], \regs[22] [0], \regs[21] [0], \regs[20] [0], 
            \regs[19] [0], \regs[18] [0], \regs[17] [0], \regs[16] [0], 
            \regs[15] [0], \regs[14] [0], \regs[13] [0], \regs[12] [0], 
            \regs[11] [0], \regs[10] [0], \regs[9] [0], \regs[8] [0], 
            \regs[7] [0], \regs[6] [0], \regs[5] [0], \regs[4] [0], 
            \regs[3] [0], \regs[2] [0], \regs[1] [0], \regs[0] [0]}), 
            .o(rd1[0]));   // regs.v(31)
    Decoder_5 Decoder_68 (.i({wa0}), .o({n69, n70, n71, n72, n73, 
            n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, 
            n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, 
            n94, n95, n96, n97, n98, n99, n100}));   // regs.v(45)
    assign n101 = n69 ? wd0[31] : pcout[31];   // regs.v(45)
    assign n102 = n69 ? wd0[30] : pcout[30];   // regs.v(45)
    assign n103 = n69 ? wd0[29] : pcout[29];   // regs.v(45)
    assign n104 = n69 ? wd0[28] : pcout[28];   // regs.v(45)
    assign n105 = n69 ? wd0[27] : pcout[27];   // regs.v(45)
    assign n106 = n69 ? wd0[26] : pcout[26];   // regs.v(45)
    assign n107 = n69 ? wd0[25] : pcout[25];   // regs.v(45)
    assign n108 = n69 ? wd0[24] : pcout[24];   // regs.v(45)
    assign n109 = n69 ? wd0[23] : pcout[23];   // regs.v(45)
    assign n110 = n69 ? wd0[22] : pcout[22];   // regs.v(45)
    assign n111 = n69 ? wd0[21] : pcout[21];   // regs.v(45)
    assign n112 = n69 ? wd0[20] : pcout[20];   // regs.v(45)
    assign n113 = n69 ? wd0[19] : pcout[19];   // regs.v(45)
    assign n114 = n69 ? wd0[18] : pcout[18];   // regs.v(45)
    assign n115 = n69 ? wd0[17] : pcout[17];   // regs.v(45)
    assign n116 = n69 ? wd0[16] : pcout[16];   // regs.v(45)
    assign n117 = n69 ? wd0[15] : pcout[15];   // regs.v(45)
    assign n118 = n69 ? wd0[14] : pcout[14];   // regs.v(45)
    assign n119 = n69 ? wd0[13] : pcout[13];   // regs.v(45)
    assign n120 = n69 ? wd0[12] : pcout[12];   // regs.v(45)
    assign n121 = n69 ? wd0[11] : pcout[11];   // regs.v(45)
    assign n122 = n69 ? wd0[10] : pcout[10];   // regs.v(45)
    assign n123 = n69 ? wd0[9] : pcout[9];   // regs.v(45)
    assign n124 = n69 ? wd0[8] : pcout[8];   // regs.v(45)
    assign n125 = n69 ? wd0[7] : pcout[7];   // regs.v(45)
    assign n126 = n69 ? wd0[6] : pcout[6];   // regs.v(45)
    assign n127 = n69 ? wd0[5] : pcout[5];   // regs.v(45)
    assign n128 = n69 ? wd0[4] : pcout[4];   // regs.v(45)
    assign n129 = n69 ? wd0[3] : pcout[3];   // regs.v(45)
    assign n130 = n69 ? wd0[2] : pcout[2];   // regs.v(45)
    assign n131 = n69 ? wd0[1] : pcout[1];   // regs.v(45)
    assign n132 = n69 ? wd0[0] : pcout[0];   // regs.v(45)
    assign n133 = n70 ? wd0[31] : spout[31];   // regs.v(45)
    assign n134 = n70 ? wd0[30] : spout[30];   // regs.v(45)
    assign n135 = n70 ? wd0[29] : spout[29];   // regs.v(45)
    assign n136 = n70 ? wd0[28] : spout[28];   // regs.v(45)
    assign n137 = n70 ? wd0[27] : spout[27];   // regs.v(45)
    assign n138 = n70 ? wd0[26] : spout[26];   // regs.v(45)
    assign n139 = n70 ? wd0[25] : spout[25];   // regs.v(45)
    assign n140 = n70 ? wd0[24] : spout[24];   // regs.v(45)
    assign n141 = n70 ? wd0[23] : spout[23];   // regs.v(45)
    assign n142 = n70 ? wd0[22] : spout[22];   // regs.v(45)
    assign n143 = n70 ? wd0[21] : spout[21];   // regs.v(45)
    assign n144 = n70 ? wd0[20] : spout[20];   // regs.v(45)
    assign n145 = n70 ? wd0[19] : spout[19];   // regs.v(45)
    assign n146 = n70 ? wd0[18] : spout[18];   // regs.v(45)
    assign n147 = n70 ? wd0[17] : spout[17];   // regs.v(45)
    assign n148 = n70 ? wd0[16] : spout[16];   // regs.v(45)
    assign n149 = n70 ? wd0[15] : spout[15];   // regs.v(45)
    assign n150 = n70 ? wd0[14] : spout[14];   // regs.v(45)
    assign n151 = n70 ? wd0[13] : spout[13];   // regs.v(45)
    assign n152 = n70 ? wd0[12] : spout[12];   // regs.v(45)
    assign n153 = n70 ? wd0[11] : spout[11];   // regs.v(45)
    assign n154 = n70 ? wd0[10] : spout[10];   // regs.v(45)
    assign n155 = n70 ? wd0[9] : spout[9];   // regs.v(45)
    assign n156 = n70 ? wd0[8] : spout[8];   // regs.v(45)
    assign n157 = n70 ? wd0[7] : spout[7];   // regs.v(45)
    assign n158 = n70 ? wd0[6] : spout[6];   // regs.v(45)
    assign n159 = n70 ? wd0[5] : spout[5];   // regs.v(45)
    assign n160 = n70 ? wd0[4] : spout[4];   // regs.v(45)
    assign n161 = n70 ? wd0[3] : spout[3];   // regs.v(45)
    assign n162 = n70 ? wd0[2] : spout[2];   // regs.v(45)
    assign n163 = n70 ? wd0[1] : spout[1];   // regs.v(45)
    assign n164 = n70 ? wd0[0] : spout[0];   // regs.v(45)
    assign n165 = n71 ? wd0[31] : lrout[31];   // regs.v(45)
    assign n166 = n71 ? wd0[30] : lrout[30];   // regs.v(45)
    assign n167 = n71 ? wd0[29] : lrout[29];   // regs.v(45)
    assign n168 = n71 ? wd0[28] : lrout[28];   // regs.v(45)
    assign n169 = n71 ? wd0[27] : lrout[27];   // regs.v(45)
    assign n170 = n71 ? wd0[26] : lrout[26];   // regs.v(45)
    assign n171 = n71 ? wd0[25] : lrout[25];   // regs.v(45)
    assign n172 = n71 ? wd0[24] : lrout[24];   // regs.v(45)
    assign n173 = n71 ? wd0[23] : lrout[23];   // regs.v(45)
    assign n174 = n71 ? wd0[22] : lrout[22];   // regs.v(45)
    assign n175 = n71 ? wd0[21] : lrout[21];   // regs.v(45)
    assign n176 = n71 ? wd0[20] : lrout[20];   // regs.v(45)
    assign n177 = n71 ? wd0[19] : lrout[19];   // regs.v(45)
    assign n178 = n71 ? wd0[18] : lrout[18];   // regs.v(45)
    assign n179 = n71 ? wd0[17] : lrout[17];   // regs.v(45)
    assign n180 = n71 ? wd0[16] : lrout[16];   // regs.v(45)
    assign n181 = n71 ? wd0[15] : lrout[15];   // regs.v(45)
    assign n182 = n71 ? wd0[14] : lrout[14];   // regs.v(45)
    assign n183 = n71 ? wd0[13] : lrout[13];   // regs.v(45)
    assign n184 = n71 ? wd0[12] : lrout[12];   // regs.v(45)
    assign n185 = n71 ? wd0[11] : lrout[11];   // regs.v(45)
    assign n186 = n71 ? wd0[10] : lrout[10];   // regs.v(45)
    assign n187 = n71 ? wd0[9] : lrout[9];   // regs.v(45)
    assign n188 = n71 ? wd0[8] : lrout[8];   // regs.v(45)
    assign n189 = n71 ? wd0[7] : lrout[7];   // regs.v(45)
    assign n190 = n71 ? wd0[6] : lrout[6];   // regs.v(45)
    assign n191 = n71 ? wd0[5] : lrout[5];   // regs.v(45)
    assign n192 = n71 ? wd0[4] : lrout[4];   // regs.v(45)
    assign n193 = n71 ? wd0[3] : lrout[3];   // regs.v(45)
    assign n194 = n71 ? wd0[2] : lrout[2];   // regs.v(45)
    assign n195 = n71 ? wd0[1] : lrout[1];   // regs.v(45)
    assign n196 = n71 ? wd0[0] : lrout[0];   // regs.v(45)
    assign n197 = n72 ? wd0[31] : stout[31];   // regs.v(45)
    assign n198 = n72 ? wd0[30] : stout[30];   // regs.v(45)
    assign n199 = n72 ? wd0[29] : stout[29];   // regs.v(45)
    assign n200 = n72 ? wd0[28] : stout[28];   // regs.v(45)
    assign n201 = n72 ? wd0[27] : stout[27];   // regs.v(45)
    assign n202 = n72 ? wd0[26] : stout[26];   // regs.v(45)
    assign n203 = n72 ? wd0[25] : stout[25];   // regs.v(45)
    assign n204 = n72 ? wd0[24] : stout[24];   // regs.v(45)
    assign n205 = n72 ? wd0[23] : stout[23];   // regs.v(45)
    assign n206 = n72 ? wd0[22] : stout[22];   // regs.v(45)
    assign n207 = n72 ? wd0[21] : stout[21];   // regs.v(45)
    assign n208 = n72 ? wd0[20] : stout[20];   // regs.v(45)
    assign n209 = n72 ? wd0[19] : stout[19];   // regs.v(45)
    assign n210 = n72 ? wd0[18] : stout[18];   // regs.v(45)
    assign n211 = n72 ? wd0[17] : stout[17];   // regs.v(45)
    assign n212 = n72 ? wd0[16] : stout[16];   // regs.v(45)
    assign n213 = n72 ? wd0[15] : stout[15];   // regs.v(45)
    assign n214 = n72 ? wd0[14] : stout[14];   // regs.v(45)
    assign n215 = n72 ? wd0[13] : stout[13];   // regs.v(45)
    assign n216 = n72 ? wd0[12] : stout[12];   // regs.v(45)
    assign n217 = n72 ? wd0[11] : stout[11];   // regs.v(45)
    assign n218 = n72 ? wd0[10] : stout[10];   // regs.v(45)
    assign n219 = n72 ? wd0[9] : stout[9];   // regs.v(45)
    assign n220 = n72 ? wd0[8] : stout[8];   // regs.v(45)
    assign n221 = n72 ? wd0[7] : stout[7];   // regs.v(45)
    assign n222 = n72 ? wd0[6] : stout[6];   // regs.v(45)
    assign n223 = n72 ? wd0[5] : stout[5];   // regs.v(45)
    assign n224 = n72 ? wd0[4] : stout[4];   // regs.v(45)
    assign n225 = n72 ? wd0[3] : stout[3];   // regs.v(45)
    assign n226 = n72 ? wd0[2] : stout[2];   // regs.v(45)
    assign n227 = n72 ? wd0[1] : stout[1];   // regs.v(45)
    assign n228 = n72 ? wd0[0] : stout[0];   // regs.v(45)
    assign n229 = n73 ? wd0[31] : \regs[27] [31];   // regs.v(45)
    assign n230 = n73 ? wd0[30] : \regs[27] [30];   // regs.v(45)
    assign n231 = n73 ? wd0[29] : \regs[27] [29];   // regs.v(45)
    assign n232 = n73 ? wd0[28] : \regs[27] [28];   // regs.v(45)
    assign n233 = n73 ? wd0[27] : \regs[27] [27];   // regs.v(45)
    assign n234 = n73 ? wd0[26] : \regs[27] [26];   // regs.v(45)
    assign n235 = n73 ? wd0[25] : \regs[27] [25];   // regs.v(45)
    assign n236 = n73 ? wd0[24] : \regs[27] [24];   // regs.v(45)
    assign n237 = n73 ? wd0[23] : \regs[27] [23];   // regs.v(45)
    assign n238 = n73 ? wd0[22] : \regs[27] [22];   // regs.v(45)
    assign n239 = n73 ? wd0[21] : \regs[27] [21];   // regs.v(45)
    assign n240 = n73 ? wd0[20] : \regs[27] [20];   // regs.v(45)
    assign n241 = n73 ? wd0[19] : \regs[27] [19];   // regs.v(45)
    assign n242 = n73 ? wd0[18] : \regs[27] [18];   // regs.v(45)
    assign n243 = n73 ? wd0[17] : \regs[27] [17];   // regs.v(45)
    assign n244 = n73 ? wd0[16] : \regs[27] [16];   // regs.v(45)
    assign n245 = n73 ? wd0[15] : \regs[27] [15];   // regs.v(45)
    assign n246 = n73 ? wd0[14] : \regs[27] [14];   // regs.v(45)
    assign n247 = n73 ? wd0[13] : \regs[27] [13];   // regs.v(45)
    assign n248 = n73 ? wd0[12] : \regs[27] [12];   // regs.v(45)
    assign n249 = n73 ? wd0[11] : \regs[27] [11];   // regs.v(45)
    assign n250 = n73 ? wd0[10] : \regs[27] [10];   // regs.v(45)
    assign n251 = n73 ? wd0[9] : \regs[27] [9];   // regs.v(45)
    assign n252 = n73 ? wd0[8] : \regs[27] [8];   // regs.v(45)
    assign n253 = n73 ? wd0[7] : \regs[27] [7];   // regs.v(45)
    assign n254 = n73 ? wd0[6] : \regs[27] [6];   // regs.v(45)
    assign n255 = n73 ? wd0[5] : \regs[27] [5];   // regs.v(45)
    assign n256 = n73 ? wd0[4] : \regs[27] [4];   // regs.v(45)
    assign n257 = n73 ? wd0[3] : \regs[27] [3];   // regs.v(45)
    assign n258 = n73 ? wd0[2] : \regs[27] [2];   // regs.v(45)
    assign n259 = n73 ? wd0[1] : \regs[27] [1];   // regs.v(45)
    assign n260 = n73 ? wd0[0] : \regs[27] [0];   // regs.v(45)
    assign n261 = n74 ? wd0[31] : \regs[26] [31];   // regs.v(45)
    assign n262 = n74 ? wd0[30] : \regs[26] [30];   // regs.v(45)
    assign n263 = n74 ? wd0[29] : \regs[26] [29];   // regs.v(45)
    assign n264 = n74 ? wd0[28] : \regs[26] [28];   // regs.v(45)
    assign n265 = n74 ? wd0[27] : \regs[26] [27];   // regs.v(45)
    assign n266 = n74 ? wd0[26] : \regs[26] [26];   // regs.v(45)
    assign n267 = n74 ? wd0[25] : \regs[26] [25];   // regs.v(45)
    assign n268 = n74 ? wd0[24] : \regs[26] [24];   // regs.v(45)
    assign n269 = n74 ? wd0[23] : \regs[26] [23];   // regs.v(45)
    assign n270 = n74 ? wd0[22] : \regs[26] [22];   // regs.v(45)
    assign n271 = n74 ? wd0[21] : \regs[26] [21];   // regs.v(45)
    assign n272 = n74 ? wd0[20] : \regs[26] [20];   // regs.v(45)
    assign n273 = n74 ? wd0[19] : \regs[26] [19];   // regs.v(45)
    assign n274 = n74 ? wd0[18] : \regs[26] [18];   // regs.v(45)
    assign n275 = n74 ? wd0[17] : \regs[26] [17];   // regs.v(45)
    assign n276 = n74 ? wd0[16] : \regs[26] [16];   // regs.v(45)
    assign n277 = n74 ? wd0[15] : \regs[26] [15];   // regs.v(45)
    assign n278 = n74 ? wd0[14] : \regs[26] [14];   // regs.v(45)
    assign n279 = n74 ? wd0[13] : \regs[26] [13];   // regs.v(45)
    assign n280 = n74 ? wd0[12] : \regs[26] [12];   // regs.v(45)
    assign n281 = n74 ? wd0[11] : \regs[26] [11];   // regs.v(45)
    assign n282 = n74 ? wd0[10] : \regs[26] [10];   // regs.v(45)
    assign n283 = n74 ? wd0[9] : \regs[26] [9];   // regs.v(45)
    assign n284 = n74 ? wd0[8] : \regs[26] [8];   // regs.v(45)
    assign n285 = n74 ? wd0[7] : \regs[26] [7];   // regs.v(45)
    assign n286 = n74 ? wd0[6] : \regs[26] [6];   // regs.v(45)
    assign n287 = n74 ? wd0[5] : \regs[26] [5];   // regs.v(45)
    assign n288 = n74 ? wd0[4] : \regs[26] [4];   // regs.v(45)
    assign n289 = n74 ? wd0[3] : \regs[26] [3];   // regs.v(45)
    assign n290 = n74 ? wd0[2] : \regs[26] [2];   // regs.v(45)
    assign n291 = n74 ? wd0[1] : \regs[26] [1];   // regs.v(45)
    assign n292 = n74 ? wd0[0] : \regs[26] [0];   // regs.v(45)
    assign n293 = n75 ? wd0[31] : \regs[25] [31];   // regs.v(45)
    assign n294 = n75 ? wd0[30] : \regs[25] [30];   // regs.v(45)
    assign n295 = n75 ? wd0[29] : \regs[25] [29];   // regs.v(45)
    assign n296 = n75 ? wd0[28] : \regs[25] [28];   // regs.v(45)
    assign n297 = n75 ? wd0[27] : \regs[25] [27];   // regs.v(45)
    assign n298 = n75 ? wd0[26] : \regs[25] [26];   // regs.v(45)
    assign n299 = n75 ? wd0[25] : \regs[25] [25];   // regs.v(45)
    assign n300 = n75 ? wd0[24] : \regs[25] [24];   // regs.v(45)
    assign n301 = n75 ? wd0[23] : \regs[25] [23];   // regs.v(45)
    assign n302 = n75 ? wd0[22] : \regs[25] [22];   // regs.v(45)
    assign n303 = n75 ? wd0[21] : \regs[25] [21];   // regs.v(45)
    assign n304 = n75 ? wd0[20] : \regs[25] [20];   // regs.v(45)
    assign n305 = n75 ? wd0[19] : \regs[25] [19];   // regs.v(45)
    assign n306 = n75 ? wd0[18] : \regs[25] [18];   // regs.v(45)
    assign n307 = n75 ? wd0[17] : \regs[25] [17];   // regs.v(45)
    assign n308 = n75 ? wd0[16] : \regs[25] [16];   // regs.v(45)
    assign n309 = n75 ? wd0[15] : \regs[25] [15];   // regs.v(45)
    assign n310 = n75 ? wd0[14] : \regs[25] [14];   // regs.v(45)
    assign n311 = n75 ? wd0[13] : \regs[25] [13];   // regs.v(45)
    assign n312 = n75 ? wd0[12] : \regs[25] [12];   // regs.v(45)
    assign n313 = n75 ? wd0[11] : \regs[25] [11];   // regs.v(45)
    assign n314 = n75 ? wd0[10] : \regs[25] [10];   // regs.v(45)
    assign n315 = n75 ? wd0[9] : \regs[25] [9];   // regs.v(45)
    assign n316 = n75 ? wd0[8] : \regs[25] [8];   // regs.v(45)
    assign n317 = n75 ? wd0[7] : \regs[25] [7];   // regs.v(45)
    assign n318 = n75 ? wd0[6] : \regs[25] [6];   // regs.v(45)
    assign n319 = n75 ? wd0[5] : \regs[25] [5];   // regs.v(45)
    assign n320 = n75 ? wd0[4] : \regs[25] [4];   // regs.v(45)
    assign n321 = n75 ? wd0[3] : \regs[25] [3];   // regs.v(45)
    assign n322 = n75 ? wd0[2] : \regs[25] [2];   // regs.v(45)
    assign n323 = n75 ? wd0[1] : \regs[25] [1];   // regs.v(45)
    assign n324 = n75 ? wd0[0] : \regs[25] [0];   // regs.v(45)
    assign n325 = n76 ? wd0[31] : \regs[24] [31];   // regs.v(45)
    assign n326 = n76 ? wd0[30] : \regs[24] [30];   // regs.v(45)
    assign n327 = n76 ? wd0[29] : \regs[24] [29];   // regs.v(45)
    assign n328 = n76 ? wd0[28] : \regs[24] [28];   // regs.v(45)
    assign n329 = n76 ? wd0[27] : \regs[24] [27];   // regs.v(45)
    assign n330 = n76 ? wd0[26] : \regs[24] [26];   // regs.v(45)
    assign n331 = n76 ? wd0[25] : \regs[24] [25];   // regs.v(45)
    assign n332 = n76 ? wd0[24] : \regs[24] [24];   // regs.v(45)
    assign n333 = n76 ? wd0[23] : \regs[24] [23];   // regs.v(45)
    assign n334 = n76 ? wd0[22] : \regs[24] [22];   // regs.v(45)
    assign n335 = n76 ? wd0[21] : \regs[24] [21];   // regs.v(45)
    assign n336 = n76 ? wd0[20] : \regs[24] [20];   // regs.v(45)
    assign n337 = n76 ? wd0[19] : \regs[24] [19];   // regs.v(45)
    assign n338 = n76 ? wd0[18] : \regs[24] [18];   // regs.v(45)
    assign n339 = n76 ? wd0[17] : \regs[24] [17];   // regs.v(45)
    assign n340 = n76 ? wd0[16] : \regs[24] [16];   // regs.v(45)
    assign n341 = n76 ? wd0[15] : \regs[24] [15];   // regs.v(45)
    assign n342 = n76 ? wd0[14] : \regs[24] [14];   // regs.v(45)
    assign n343 = n76 ? wd0[13] : \regs[24] [13];   // regs.v(45)
    assign n344 = n76 ? wd0[12] : \regs[24] [12];   // regs.v(45)
    assign n345 = n76 ? wd0[11] : \regs[24] [11];   // regs.v(45)
    assign n346 = n76 ? wd0[10] : \regs[24] [10];   // regs.v(45)
    assign n347 = n76 ? wd0[9] : \regs[24] [9];   // regs.v(45)
    assign n348 = n76 ? wd0[8] : \regs[24] [8];   // regs.v(45)
    assign n349 = n76 ? wd0[7] : \regs[24] [7];   // regs.v(45)
    assign n350 = n76 ? wd0[6] : \regs[24] [6];   // regs.v(45)
    assign n351 = n76 ? wd0[5] : \regs[24] [5];   // regs.v(45)
    assign n352 = n76 ? wd0[4] : \regs[24] [4];   // regs.v(45)
    assign n353 = n76 ? wd0[3] : \regs[24] [3];   // regs.v(45)
    assign n354 = n76 ? wd0[2] : \regs[24] [2];   // regs.v(45)
    assign n355 = n76 ? wd0[1] : \regs[24] [1];   // regs.v(45)
    assign n356 = n76 ? wd0[0] : \regs[24] [0];   // regs.v(45)
    assign n357 = n77 ? wd0[31] : \regs[23] [31];   // regs.v(45)
    assign n358 = n77 ? wd0[30] : \regs[23] [30];   // regs.v(45)
    assign n359 = n77 ? wd0[29] : \regs[23] [29];   // regs.v(45)
    assign n360 = n77 ? wd0[28] : \regs[23] [28];   // regs.v(45)
    assign n361 = n77 ? wd0[27] : \regs[23] [27];   // regs.v(45)
    assign n362 = n77 ? wd0[26] : \regs[23] [26];   // regs.v(45)
    assign n363 = n77 ? wd0[25] : \regs[23] [25];   // regs.v(45)
    assign n364 = n77 ? wd0[24] : \regs[23] [24];   // regs.v(45)
    assign n365 = n77 ? wd0[23] : \regs[23] [23];   // regs.v(45)
    assign n366 = n77 ? wd0[22] : \regs[23] [22];   // regs.v(45)
    assign n367 = n77 ? wd0[21] : \regs[23] [21];   // regs.v(45)
    assign n368 = n77 ? wd0[20] : \regs[23] [20];   // regs.v(45)
    assign n369 = n77 ? wd0[19] : \regs[23] [19];   // regs.v(45)
    assign n370 = n77 ? wd0[18] : \regs[23] [18];   // regs.v(45)
    assign n371 = n77 ? wd0[17] : \regs[23] [17];   // regs.v(45)
    assign n372 = n77 ? wd0[16] : \regs[23] [16];   // regs.v(45)
    assign n373 = n77 ? wd0[15] : \regs[23] [15];   // regs.v(45)
    assign n374 = n77 ? wd0[14] : \regs[23] [14];   // regs.v(45)
    assign n375 = n77 ? wd0[13] : \regs[23] [13];   // regs.v(45)
    assign n376 = n77 ? wd0[12] : \regs[23] [12];   // regs.v(45)
    assign n377 = n77 ? wd0[11] : \regs[23] [11];   // regs.v(45)
    assign n378 = n77 ? wd0[10] : \regs[23] [10];   // regs.v(45)
    assign n379 = n77 ? wd0[9] : \regs[23] [9];   // regs.v(45)
    assign n380 = n77 ? wd0[8] : \regs[23] [8];   // regs.v(45)
    assign n381 = n77 ? wd0[7] : \regs[23] [7];   // regs.v(45)
    assign n382 = n77 ? wd0[6] : \regs[23] [6];   // regs.v(45)
    assign n383 = n77 ? wd0[5] : \regs[23] [5];   // regs.v(45)
    assign n384 = n77 ? wd0[4] : \regs[23] [4];   // regs.v(45)
    assign n385 = n77 ? wd0[3] : \regs[23] [3];   // regs.v(45)
    assign n386 = n77 ? wd0[2] : \regs[23] [2];   // regs.v(45)
    assign n387 = n77 ? wd0[1] : \regs[23] [1];   // regs.v(45)
    assign n388 = n77 ? wd0[0] : \regs[23] [0];   // regs.v(45)
    assign n389 = n78 ? wd0[31] : \regs[22] [31];   // regs.v(45)
    assign n390 = n78 ? wd0[30] : \regs[22] [30];   // regs.v(45)
    assign n391 = n78 ? wd0[29] : \regs[22] [29];   // regs.v(45)
    assign n392 = n78 ? wd0[28] : \regs[22] [28];   // regs.v(45)
    assign n393 = n78 ? wd0[27] : \regs[22] [27];   // regs.v(45)
    assign n394 = n78 ? wd0[26] : \regs[22] [26];   // regs.v(45)
    assign n395 = n78 ? wd0[25] : \regs[22] [25];   // regs.v(45)
    assign n396 = n78 ? wd0[24] : \regs[22] [24];   // regs.v(45)
    assign n397 = n78 ? wd0[23] : \regs[22] [23];   // regs.v(45)
    assign n398 = n78 ? wd0[22] : \regs[22] [22];   // regs.v(45)
    assign n399 = n78 ? wd0[21] : \regs[22] [21];   // regs.v(45)
    assign n400 = n78 ? wd0[20] : \regs[22] [20];   // regs.v(45)
    assign n401 = n78 ? wd0[19] : \regs[22] [19];   // regs.v(45)
    assign n402 = n78 ? wd0[18] : \regs[22] [18];   // regs.v(45)
    assign n403 = n78 ? wd0[17] : \regs[22] [17];   // regs.v(45)
    assign n404 = n78 ? wd0[16] : \regs[22] [16];   // regs.v(45)
    assign n405 = n78 ? wd0[15] : \regs[22] [15];   // regs.v(45)
    assign n406 = n78 ? wd0[14] : \regs[22] [14];   // regs.v(45)
    assign n407 = n78 ? wd0[13] : \regs[22] [13];   // regs.v(45)
    assign n408 = n78 ? wd0[12] : \regs[22] [12];   // regs.v(45)
    assign n409 = n78 ? wd0[11] : \regs[22] [11];   // regs.v(45)
    assign n410 = n78 ? wd0[10] : \regs[22] [10];   // regs.v(45)
    assign n411 = n78 ? wd0[9] : \regs[22] [9];   // regs.v(45)
    assign n412 = n78 ? wd0[8] : \regs[22] [8];   // regs.v(45)
    assign n413 = n78 ? wd0[7] : \regs[22] [7];   // regs.v(45)
    assign n414 = n78 ? wd0[6] : \regs[22] [6];   // regs.v(45)
    assign n415 = n78 ? wd0[5] : \regs[22] [5];   // regs.v(45)
    assign n416 = n78 ? wd0[4] : \regs[22] [4];   // regs.v(45)
    assign n417 = n78 ? wd0[3] : \regs[22] [3];   // regs.v(45)
    assign n418 = n78 ? wd0[2] : \regs[22] [2];   // regs.v(45)
    assign n419 = n78 ? wd0[1] : \regs[22] [1];   // regs.v(45)
    assign n420 = n78 ? wd0[0] : \regs[22] [0];   // regs.v(45)
    assign n421 = n79 ? wd0[31] : \regs[21] [31];   // regs.v(45)
    assign n422 = n79 ? wd0[30] : \regs[21] [30];   // regs.v(45)
    assign n423 = n79 ? wd0[29] : \regs[21] [29];   // regs.v(45)
    assign n424 = n79 ? wd0[28] : \regs[21] [28];   // regs.v(45)
    assign n425 = n79 ? wd0[27] : \regs[21] [27];   // regs.v(45)
    assign n426 = n79 ? wd0[26] : \regs[21] [26];   // regs.v(45)
    assign n427 = n79 ? wd0[25] : \regs[21] [25];   // regs.v(45)
    assign n428 = n79 ? wd0[24] : \regs[21] [24];   // regs.v(45)
    assign n429 = n79 ? wd0[23] : \regs[21] [23];   // regs.v(45)
    assign n430 = n79 ? wd0[22] : \regs[21] [22];   // regs.v(45)
    assign n431 = n79 ? wd0[21] : \regs[21] [21];   // regs.v(45)
    assign n432 = n79 ? wd0[20] : \regs[21] [20];   // regs.v(45)
    assign n433 = n79 ? wd0[19] : \regs[21] [19];   // regs.v(45)
    assign n434 = n79 ? wd0[18] : \regs[21] [18];   // regs.v(45)
    assign n435 = n79 ? wd0[17] : \regs[21] [17];   // regs.v(45)
    assign n436 = n79 ? wd0[16] : \regs[21] [16];   // regs.v(45)
    assign n437 = n79 ? wd0[15] : \regs[21] [15];   // regs.v(45)
    assign n438 = n79 ? wd0[14] : \regs[21] [14];   // regs.v(45)
    assign n439 = n79 ? wd0[13] : \regs[21] [13];   // regs.v(45)
    assign n440 = n79 ? wd0[12] : \regs[21] [12];   // regs.v(45)
    assign n441 = n79 ? wd0[11] : \regs[21] [11];   // regs.v(45)
    assign n442 = n79 ? wd0[10] : \regs[21] [10];   // regs.v(45)
    assign n443 = n79 ? wd0[9] : \regs[21] [9];   // regs.v(45)
    assign n444 = n79 ? wd0[8] : \regs[21] [8];   // regs.v(45)
    assign n445 = n79 ? wd0[7] : \regs[21] [7];   // regs.v(45)
    assign n446 = n79 ? wd0[6] : \regs[21] [6];   // regs.v(45)
    assign n447 = n79 ? wd0[5] : \regs[21] [5];   // regs.v(45)
    assign n448 = n79 ? wd0[4] : \regs[21] [4];   // regs.v(45)
    assign n449 = n79 ? wd0[3] : \regs[21] [3];   // regs.v(45)
    assign n450 = n79 ? wd0[2] : \regs[21] [2];   // regs.v(45)
    assign n451 = n79 ? wd0[1] : \regs[21] [1];   // regs.v(45)
    assign n452 = n79 ? wd0[0] : \regs[21] [0];   // regs.v(45)
    assign n453 = n80 ? wd0[31] : \regs[20] [31];   // regs.v(45)
    assign n454 = n80 ? wd0[30] : \regs[20] [30];   // regs.v(45)
    assign n455 = n80 ? wd0[29] : \regs[20] [29];   // regs.v(45)
    assign n456 = n80 ? wd0[28] : \regs[20] [28];   // regs.v(45)
    assign n457 = n80 ? wd0[27] : \regs[20] [27];   // regs.v(45)
    assign n458 = n80 ? wd0[26] : \regs[20] [26];   // regs.v(45)
    assign n459 = n80 ? wd0[25] : \regs[20] [25];   // regs.v(45)
    assign n460 = n80 ? wd0[24] : \regs[20] [24];   // regs.v(45)
    assign n461 = n80 ? wd0[23] : \regs[20] [23];   // regs.v(45)
    assign n462 = n80 ? wd0[22] : \regs[20] [22];   // regs.v(45)
    assign n463 = n80 ? wd0[21] : \regs[20] [21];   // regs.v(45)
    assign n464 = n80 ? wd0[20] : \regs[20] [20];   // regs.v(45)
    assign n465 = n80 ? wd0[19] : \regs[20] [19];   // regs.v(45)
    assign n466 = n80 ? wd0[18] : \regs[20] [18];   // regs.v(45)
    assign n467 = n80 ? wd0[17] : \regs[20] [17];   // regs.v(45)
    assign n468 = n80 ? wd0[16] : \regs[20] [16];   // regs.v(45)
    assign n469 = n80 ? wd0[15] : \regs[20] [15];   // regs.v(45)
    assign n470 = n80 ? wd0[14] : \regs[20] [14];   // regs.v(45)
    assign n471 = n80 ? wd0[13] : \regs[20] [13];   // regs.v(45)
    assign n472 = n80 ? wd0[12] : \regs[20] [12];   // regs.v(45)
    assign n473 = n80 ? wd0[11] : \regs[20] [11];   // regs.v(45)
    assign n474 = n80 ? wd0[10] : \regs[20] [10];   // regs.v(45)
    assign n475 = n80 ? wd0[9] : \regs[20] [9];   // regs.v(45)
    assign n476 = n80 ? wd0[8] : \regs[20] [8];   // regs.v(45)
    assign n477 = n80 ? wd0[7] : \regs[20] [7];   // regs.v(45)
    assign n478 = n80 ? wd0[6] : \regs[20] [6];   // regs.v(45)
    assign n479 = n80 ? wd0[5] : \regs[20] [5];   // regs.v(45)
    assign n480 = n80 ? wd0[4] : \regs[20] [4];   // regs.v(45)
    assign n481 = n80 ? wd0[3] : \regs[20] [3];   // regs.v(45)
    assign n482 = n80 ? wd0[2] : \regs[20] [2];   // regs.v(45)
    assign n483 = n80 ? wd0[1] : \regs[20] [1];   // regs.v(45)
    assign n484 = n80 ? wd0[0] : \regs[20] [0];   // regs.v(45)
    assign n485 = n81 ? wd0[31] : \regs[19] [31];   // regs.v(45)
    assign n486 = n81 ? wd0[30] : \regs[19] [30];   // regs.v(45)
    assign n487 = n81 ? wd0[29] : \regs[19] [29];   // regs.v(45)
    assign n488 = n81 ? wd0[28] : \regs[19] [28];   // regs.v(45)
    assign n489 = n81 ? wd0[27] : \regs[19] [27];   // regs.v(45)
    assign n490 = n81 ? wd0[26] : \regs[19] [26];   // regs.v(45)
    assign n491 = n81 ? wd0[25] : \regs[19] [25];   // regs.v(45)
    assign n492 = n81 ? wd0[24] : \regs[19] [24];   // regs.v(45)
    assign n493 = n81 ? wd0[23] : \regs[19] [23];   // regs.v(45)
    assign n494 = n81 ? wd0[22] : \regs[19] [22];   // regs.v(45)
    assign n495 = n81 ? wd0[21] : \regs[19] [21];   // regs.v(45)
    assign n496 = n81 ? wd0[20] : \regs[19] [20];   // regs.v(45)
    assign n497 = n81 ? wd0[19] : \regs[19] [19];   // regs.v(45)
    assign n498 = n81 ? wd0[18] : \regs[19] [18];   // regs.v(45)
    assign n499 = n81 ? wd0[17] : \regs[19] [17];   // regs.v(45)
    assign n500 = n81 ? wd0[16] : \regs[19] [16];   // regs.v(45)
    assign n501 = n81 ? wd0[15] : \regs[19] [15];   // regs.v(45)
    assign n502 = n81 ? wd0[14] : \regs[19] [14];   // regs.v(45)
    assign n503 = n81 ? wd0[13] : \regs[19] [13];   // regs.v(45)
    assign n504 = n81 ? wd0[12] : \regs[19] [12];   // regs.v(45)
    assign n505 = n81 ? wd0[11] : \regs[19] [11];   // regs.v(45)
    assign n506 = n81 ? wd0[10] : \regs[19] [10];   // regs.v(45)
    assign n507 = n81 ? wd0[9] : \regs[19] [9];   // regs.v(45)
    assign n508 = n81 ? wd0[8] : \regs[19] [8];   // regs.v(45)
    assign n509 = n81 ? wd0[7] : \regs[19] [7];   // regs.v(45)
    assign n510 = n81 ? wd0[6] : \regs[19] [6];   // regs.v(45)
    assign n511 = n81 ? wd0[5] : \regs[19] [5];   // regs.v(45)
    assign n512 = n81 ? wd0[4] : \regs[19] [4];   // regs.v(45)
    assign n513 = n81 ? wd0[3] : \regs[19] [3];   // regs.v(45)
    assign n514 = n81 ? wd0[2] : \regs[19] [2];   // regs.v(45)
    assign n515 = n81 ? wd0[1] : \regs[19] [1];   // regs.v(45)
    assign n516 = n81 ? wd0[0] : \regs[19] [0];   // regs.v(45)
    assign n517 = n82 ? wd0[31] : \regs[18] [31];   // regs.v(45)
    assign n518 = n82 ? wd0[30] : \regs[18] [30];   // regs.v(45)
    assign n519 = n82 ? wd0[29] : \regs[18] [29];   // regs.v(45)
    assign n520 = n82 ? wd0[28] : \regs[18] [28];   // regs.v(45)
    assign n521 = n82 ? wd0[27] : \regs[18] [27];   // regs.v(45)
    assign n522 = n82 ? wd0[26] : \regs[18] [26];   // regs.v(45)
    assign n523 = n82 ? wd0[25] : \regs[18] [25];   // regs.v(45)
    assign n524 = n82 ? wd0[24] : \regs[18] [24];   // regs.v(45)
    assign n525 = n82 ? wd0[23] : \regs[18] [23];   // regs.v(45)
    assign n526 = n82 ? wd0[22] : \regs[18] [22];   // regs.v(45)
    assign n527 = n82 ? wd0[21] : \regs[18] [21];   // regs.v(45)
    assign n528 = n82 ? wd0[20] : \regs[18] [20];   // regs.v(45)
    assign n529 = n82 ? wd0[19] : \regs[18] [19];   // regs.v(45)
    assign n530 = n82 ? wd0[18] : \regs[18] [18];   // regs.v(45)
    assign n531 = n82 ? wd0[17] : \regs[18] [17];   // regs.v(45)
    assign n532 = n82 ? wd0[16] : \regs[18] [16];   // regs.v(45)
    assign n533 = n82 ? wd0[15] : \regs[18] [15];   // regs.v(45)
    assign n534 = n82 ? wd0[14] : \regs[18] [14];   // regs.v(45)
    assign n535 = n82 ? wd0[13] : \regs[18] [13];   // regs.v(45)
    assign n536 = n82 ? wd0[12] : \regs[18] [12];   // regs.v(45)
    assign n537 = n82 ? wd0[11] : \regs[18] [11];   // regs.v(45)
    assign n538 = n82 ? wd0[10] : \regs[18] [10];   // regs.v(45)
    assign n539 = n82 ? wd0[9] : \regs[18] [9];   // regs.v(45)
    assign n540 = n82 ? wd0[8] : \regs[18] [8];   // regs.v(45)
    assign n541 = n82 ? wd0[7] : \regs[18] [7];   // regs.v(45)
    assign n542 = n82 ? wd0[6] : \regs[18] [6];   // regs.v(45)
    assign n543 = n82 ? wd0[5] : \regs[18] [5];   // regs.v(45)
    assign n544 = n82 ? wd0[4] : \regs[18] [4];   // regs.v(45)
    assign n545 = n82 ? wd0[3] : \regs[18] [3];   // regs.v(45)
    assign n546 = n82 ? wd0[2] : \regs[18] [2];   // regs.v(45)
    assign n547 = n82 ? wd0[1] : \regs[18] [1];   // regs.v(45)
    assign n548 = n82 ? wd0[0] : \regs[18] [0];   // regs.v(45)
    assign n549 = n83 ? wd0[31] : \regs[17] [31];   // regs.v(45)
    assign n550 = n83 ? wd0[30] : \regs[17] [30];   // regs.v(45)
    assign n551 = n83 ? wd0[29] : \regs[17] [29];   // regs.v(45)
    assign n552 = n83 ? wd0[28] : \regs[17] [28];   // regs.v(45)
    assign n553 = n83 ? wd0[27] : \regs[17] [27];   // regs.v(45)
    assign n554 = n83 ? wd0[26] : \regs[17] [26];   // regs.v(45)
    assign n555 = n83 ? wd0[25] : \regs[17] [25];   // regs.v(45)
    assign n556 = n83 ? wd0[24] : \regs[17] [24];   // regs.v(45)
    assign n557 = n83 ? wd0[23] : \regs[17] [23];   // regs.v(45)
    assign n558 = n83 ? wd0[22] : \regs[17] [22];   // regs.v(45)
    assign n559 = n83 ? wd0[21] : \regs[17] [21];   // regs.v(45)
    assign n560 = n83 ? wd0[20] : \regs[17] [20];   // regs.v(45)
    assign n561 = n83 ? wd0[19] : \regs[17] [19];   // regs.v(45)
    assign n562 = n83 ? wd0[18] : \regs[17] [18];   // regs.v(45)
    assign n563 = n83 ? wd0[17] : \regs[17] [17];   // regs.v(45)
    assign n564 = n83 ? wd0[16] : \regs[17] [16];   // regs.v(45)
    assign n565 = n83 ? wd0[15] : \regs[17] [15];   // regs.v(45)
    assign n566 = n83 ? wd0[14] : \regs[17] [14];   // regs.v(45)
    assign n567 = n83 ? wd0[13] : \regs[17] [13];   // regs.v(45)
    assign n568 = n83 ? wd0[12] : \regs[17] [12];   // regs.v(45)
    assign n569 = n83 ? wd0[11] : \regs[17] [11];   // regs.v(45)
    assign n570 = n83 ? wd0[10] : \regs[17] [10];   // regs.v(45)
    assign n571 = n83 ? wd0[9] : \regs[17] [9];   // regs.v(45)
    assign n572 = n83 ? wd0[8] : \regs[17] [8];   // regs.v(45)
    assign n573 = n83 ? wd0[7] : \regs[17] [7];   // regs.v(45)
    assign n574 = n83 ? wd0[6] : \regs[17] [6];   // regs.v(45)
    assign n575 = n83 ? wd0[5] : \regs[17] [5];   // regs.v(45)
    assign n576 = n83 ? wd0[4] : \regs[17] [4];   // regs.v(45)
    assign n577 = n83 ? wd0[3] : \regs[17] [3];   // regs.v(45)
    assign n578 = n83 ? wd0[2] : \regs[17] [2];   // regs.v(45)
    assign n579 = n83 ? wd0[1] : \regs[17] [1];   // regs.v(45)
    assign n580 = n83 ? wd0[0] : \regs[17] [0];   // regs.v(45)
    assign n581 = n84 ? wd0[31] : \regs[16] [31];   // regs.v(45)
    assign n582 = n84 ? wd0[30] : \regs[16] [30];   // regs.v(45)
    assign n583 = n84 ? wd0[29] : \regs[16] [29];   // regs.v(45)
    assign n584 = n84 ? wd0[28] : \regs[16] [28];   // regs.v(45)
    assign n585 = n84 ? wd0[27] : \regs[16] [27];   // regs.v(45)
    assign n586 = n84 ? wd0[26] : \regs[16] [26];   // regs.v(45)
    assign n587 = n84 ? wd0[25] : \regs[16] [25];   // regs.v(45)
    assign n588 = n84 ? wd0[24] : \regs[16] [24];   // regs.v(45)
    assign n589 = n84 ? wd0[23] : \regs[16] [23];   // regs.v(45)
    assign n590 = n84 ? wd0[22] : \regs[16] [22];   // regs.v(45)
    assign n591 = n84 ? wd0[21] : \regs[16] [21];   // regs.v(45)
    assign n592 = n84 ? wd0[20] : \regs[16] [20];   // regs.v(45)
    assign n593 = n84 ? wd0[19] : \regs[16] [19];   // regs.v(45)
    assign n594 = n84 ? wd0[18] : \regs[16] [18];   // regs.v(45)
    assign n595 = n84 ? wd0[17] : \regs[16] [17];   // regs.v(45)
    assign n596 = n84 ? wd0[16] : \regs[16] [16];   // regs.v(45)
    assign n597 = n84 ? wd0[15] : \regs[16] [15];   // regs.v(45)
    assign n598 = n84 ? wd0[14] : \regs[16] [14];   // regs.v(45)
    assign n599 = n84 ? wd0[13] : \regs[16] [13];   // regs.v(45)
    assign n600 = n84 ? wd0[12] : \regs[16] [12];   // regs.v(45)
    assign n601 = n84 ? wd0[11] : \regs[16] [11];   // regs.v(45)
    assign n602 = n84 ? wd0[10] : \regs[16] [10];   // regs.v(45)
    assign n603 = n84 ? wd0[9] : \regs[16] [9];   // regs.v(45)
    assign n604 = n84 ? wd0[8] : \regs[16] [8];   // regs.v(45)
    assign n605 = n84 ? wd0[7] : \regs[16] [7];   // regs.v(45)
    assign n606 = n84 ? wd0[6] : \regs[16] [6];   // regs.v(45)
    assign n607 = n84 ? wd0[5] : \regs[16] [5];   // regs.v(45)
    assign n608 = n84 ? wd0[4] : \regs[16] [4];   // regs.v(45)
    assign n609 = n84 ? wd0[3] : \regs[16] [3];   // regs.v(45)
    assign n610 = n84 ? wd0[2] : \regs[16] [2];   // regs.v(45)
    assign n611 = n84 ? wd0[1] : \regs[16] [1];   // regs.v(45)
    assign n612 = n84 ? wd0[0] : \regs[16] [0];   // regs.v(45)
    assign n613 = n85 ? wd0[31] : \regs[15] [31];   // regs.v(45)
    assign n614 = n85 ? wd0[30] : \regs[15] [30];   // regs.v(45)
    assign n615 = n85 ? wd0[29] : \regs[15] [29];   // regs.v(45)
    assign n616 = n85 ? wd0[28] : \regs[15] [28];   // regs.v(45)
    assign n617 = n85 ? wd0[27] : \regs[15] [27];   // regs.v(45)
    assign n618 = n85 ? wd0[26] : \regs[15] [26];   // regs.v(45)
    assign n619 = n85 ? wd0[25] : \regs[15] [25];   // regs.v(45)
    assign n620 = n85 ? wd0[24] : \regs[15] [24];   // regs.v(45)
    assign n621 = n85 ? wd0[23] : \regs[15] [23];   // regs.v(45)
    assign n622 = n85 ? wd0[22] : \regs[15] [22];   // regs.v(45)
    assign n623 = n85 ? wd0[21] : \regs[15] [21];   // regs.v(45)
    assign n624 = n85 ? wd0[20] : \regs[15] [20];   // regs.v(45)
    assign n625 = n85 ? wd0[19] : \regs[15] [19];   // regs.v(45)
    assign n626 = n85 ? wd0[18] : \regs[15] [18];   // regs.v(45)
    assign n627 = n85 ? wd0[17] : \regs[15] [17];   // regs.v(45)
    assign n628 = n85 ? wd0[16] : \regs[15] [16];   // regs.v(45)
    assign n629 = n85 ? wd0[15] : \regs[15] [15];   // regs.v(45)
    assign n630 = n85 ? wd0[14] : \regs[15] [14];   // regs.v(45)
    assign n631 = n85 ? wd0[13] : \regs[15] [13];   // regs.v(45)
    assign n632 = n85 ? wd0[12] : \regs[15] [12];   // regs.v(45)
    assign n633 = n85 ? wd0[11] : \regs[15] [11];   // regs.v(45)
    assign n634 = n85 ? wd0[10] : \regs[15] [10];   // regs.v(45)
    assign n635 = n85 ? wd0[9] : \regs[15] [9];   // regs.v(45)
    assign n636 = n85 ? wd0[8] : \regs[15] [8];   // regs.v(45)
    assign n637 = n85 ? wd0[7] : \regs[15] [7];   // regs.v(45)
    assign n638 = n85 ? wd0[6] : \regs[15] [6];   // regs.v(45)
    assign n639 = n85 ? wd0[5] : \regs[15] [5];   // regs.v(45)
    assign n640 = n85 ? wd0[4] : \regs[15] [4];   // regs.v(45)
    assign n641 = n85 ? wd0[3] : \regs[15] [3];   // regs.v(45)
    assign n642 = n85 ? wd0[2] : \regs[15] [2];   // regs.v(45)
    assign n643 = n85 ? wd0[1] : \regs[15] [1];   // regs.v(45)
    assign n644 = n85 ? wd0[0] : \regs[15] [0];   // regs.v(45)
    assign n645 = n86 ? wd0[31] : \regs[14] [31];   // regs.v(45)
    assign n646 = n86 ? wd0[30] : \regs[14] [30];   // regs.v(45)
    assign n647 = n86 ? wd0[29] : \regs[14] [29];   // regs.v(45)
    assign n648 = n86 ? wd0[28] : \regs[14] [28];   // regs.v(45)
    assign n649 = n86 ? wd0[27] : \regs[14] [27];   // regs.v(45)
    assign n650 = n86 ? wd0[26] : \regs[14] [26];   // regs.v(45)
    assign n651 = n86 ? wd0[25] : \regs[14] [25];   // regs.v(45)
    assign n652 = n86 ? wd0[24] : \regs[14] [24];   // regs.v(45)
    assign n653 = n86 ? wd0[23] : \regs[14] [23];   // regs.v(45)
    assign n654 = n86 ? wd0[22] : \regs[14] [22];   // regs.v(45)
    assign n655 = n86 ? wd0[21] : \regs[14] [21];   // regs.v(45)
    assign n656 = n86 ? wd0[20] : \regs[14] [20];   // regs.v(45)
    assign n657 = n86 ? wd0[19] : \regs[14] [19];   // regs.v(45)
    assign n658 = n86 ? wd0[18] : \regs[14] [18];   // regs.v(45)
    assign n659 = n86 ? wd0[17] : \regs[14] [17];   // regs.v(45)
    assign n660 = n86 ? wd0[16] : \regs[14] [16];   // regs.v(45)
    assign n661 = n86 ? wd0[15] : \regs[14] [15];   // regs.v(45)
    assign n662 = n86 ? wd0[14] : \regs[14] [14];   // regs.v(45)
    assign n663 = n86 ? wd0[13] : \regs[14] [13];   // regs.v(45)
    assign n664 = n86 ? wd0[12] : \regs[14] [12];   // regs.v(45)
    assign n665 = n86 ? wd0[11] : \regs[14] [11];   // regs.v(45)
    assign n666 = n86 ? wd0[10] : \regs[14] [10];   // regs.v(45)
    assign n667 = n86 ? wd0[9] : \regs[14] [9];   // regs.v(45)
    assign n668 = n86 ? wd0[8] : \regs[14] [8];   // regs.v(45)
    assign n669 = n86 ? wd0[7] : \regs[14] [7];   // regs.v(45)
    assign n670 = n86 ? wd0[6] : \regs[14] [6];   // regs.v(45)
    assign n671 = n86 ? wd0[5] : \regs[14] [5];   // regs.v(45)
    assign n672 = n86 ? wd0[4] : \regs[14] [4];   // regs.v(45)
    assign n673 = n86 ? wd0[3] : \regs[14] [3];   // regs.v(45)
    assign n674 = n86 ? wd0[2] : \regs[14] [2];   // regs.v(45)
    assign n675 = n86 ? wd0[1] : \regs[14] [1];   // regs.v(45)
    assign n676 = n86 ? wd0[0] : \regs[14] [0];   // regs.v(45)
    assign n677 = n87 ? wd0[31] : \regs[13] [31];   // regs.v(45)
    assign n678 = n87 ? wd0[30] : \regs[13] [30];   // regs.v(45)
    assign n679 = n87 ? wd0[29] : \regs[13] [29];   // regs.v(45)
    assign n680 = n87 ? wd0[28] : \regs[13] [28];   // regs.v(45)
    assign n681 = n87 ? wd0[27] : \regs[13] [27];   // regs.v(45)
    assign n682 = n87 ? wd0[26] : \regs[13] [26];   // regs.v(45)
    assign n683 = n87 ? wd0[25] : \regs[13] [25];   // regs.v(45)
    assign n684 = n87 ? wd0[24] : \regs[13] [24];   // regs.v(45)
    assign n685 = n87 ? wd0[23] : \regs[13] [23];   // regs.v(45)
    assign n686 = n87 ? wd0[22] : \regs[13] [22];   // regs.v(45)
    assign n687 = n87 ? wd0[21] : \regs[13] [21];   // regs.v(45)
    assign n688 = n87 ? wd0[20] : \regs[13] [20];   // regs.v(45)
    assign n689 = n87 ? wd0[19] : \regs[13] [19];   // regs.v(45)
    assign n690 = n87 ? wd0[18] : \regs[13] [18];   // regs.v(45)
    assign n691 = n87 ? wd0[17] : \regs[13] [17];   // regs.v(45)
    assign n692 = n87 ? wd0[16] : \regs[13] [16];   // regs.v(45)
    assign n693 = n87 ? wd0[15] : \regs[13] [15];   // regs.v(45)
    assign n694 = n87 ? wd0[14] : \regs[13] [14];   // regs.v(45)
    assign n695 = n87 ? wd0[13] : \regs[13] [13];   // regs.v(45)
    assign n696 = n87 ? wd0[12] : \regs[13] [12];   // regs.v(45)
    assign n697 = n87 ? wd0[11] : \regs[13] [11];   // regs.v(45)
    assign n698 = n87 ? wd0[10] : \regs[13] [10];   // regs.v(45)
    assign n699 = n87 ? wd0[9] : \regs[13] [9];   // regs.v(45)
    assign n700 = n87 ? wd0[8] : \regs[13] [8];   // regs.v(45)
    assign n701 = n87 ? wd0[7] : \regs[13] [7];   // regs.v(45)
    assign n702 = n87 ? wd0[6] : \regs[13] [6];   // regs.v(45)
    assign n703 = n87 ? wd0[5] : \regs[13] [5];   // regs.v(45)
    assign n704 = n87 ? wd0[4] : \regs[13] [4];   // regs.v(45)
    assign n705 = n87 ? wd0[3] : \regs[13] [3];   // regs.v(45)
    assign n706 = n87 ? wd0[2] : \regs[13] [2];   // regs.v(45)
    assign n707 = n87 ? wd0[1] : \regs[13] [1];   // regs.v(45)
    assign n708 = n87 ? wd0[0] : \regs[13] [0];   // regs.v(45)
    assign n709 = n88 ? wd0[31] : \regs[12] [31];   // regs.v(45)
    assign n710 = n88 ? wd0[30] : \regs[12] [30];   // regs.v(45)
    assign n711 = n88 ? wd0[29] : \regs[12] [29];   // regs.v(45)
    assign n712 = n88 ? wd0[28] : \regs[12] [28];   // regs.v(45)
    assign n713 = n88 ? wd0[27] : \regs[12] [27];   // regs.v(45)
    assign n714 = n88 ? wd0[26] : \regs[12] [26];   // regs.v(45)
    assign n715 = n88 ? wd0[25] : \regs[12] [25];   // regs.v(45)
    assign n716 = n88 ? wd0[24] : \regs[12] [24];   // regs.v(45)
    assign n717 = n88 ? wd0[23] : \regs[12] [23];   // regs.v(45)
    assign n718 = n88 ? wd0[22] : \regs[12] [22];   // regs.v(45)
    assign n719 = n88 ? wd0[21] : \regs[12] [21];   // regs.v(45)
    assign n720 = n88 ? wd0[20] : \regs[12] [20];   // regs.v(45)
    assign n721 = n88 ? wd0[19] : \regs[12] [19];   // regs.v(45)
    assign n722 = n88 ? wd0[18] : \regs[12] [18];   // regs.v(45)
    assign n723 = n88 ? wd0[17] : \regs[12] [17];   // regs.v(45)
    assign n724 = n88 ? wd0[16] : \regs[12] [16];   // regs.v(45)
    assign n725 = n88 ? wd0[15] : \regs[12] [15];   // regs.v(45)
    assign n726 = n88 ? wd0[14] : \regs[12] [14];   // regs.v(45)
    assign n727 = n88 ? wd0[13] : \regs[12] [13];   // regs.v(45)
    assign n728 = n88 ? wd0[12] : \regs[12] [12];   // regs.v(45)
    assign n729 = n88 ? wd0[11] : \regs[12] [11];   // regs.v(45)
    assign n730 = n88 ? wd0[10] : \regs[12] [10];   // regs.v(45)
    assign n731 = n88 ? wd0[9] : \regs[12] [9];   // regs.v(45)
    assign n732 = n88 ? wd0[8] : \regs[12] [8];   // regs.v(45)
    assign n733 = n88 ? wd0[7] : \regs[12] [7];   // regs.v(45)
    assign n734 = n88 ? wd0[6] : \regs[12] [6];   // regs.v(45)
    assign n735 = n88 ? wd0[5] : \regs[12] [5];   // regs.v(45)
    assign n736 = n88 ? wd0[4] : \regs[12] [4];   // regs.v(45)
    assign n737 = n88 ? wd0[3] : \regs[12] [3];   // regs.v(45)
    assign n738 = n88 ? wd0[2] : \regs[12] [2];   // regs.v(45)
    assign n739 = n88 ? wd0[1] : \regs[12] [1];   // regs.v(45)
    assign n740 = n88 ? wd0[0] : \regs[12] [0];   // regs.v(45)
    assign n741 = n89 ? wd0[31] : \regs[11] [31];   // regs.v(45)
    assign n742 = n89 ? wd0[30] : \regs[11] [30];   // regs.v(45)
    assign n743 = n89 ? wd0[29] : \regs[11] [29];   // regs.v(45)
    assign n744 = n89 ? wd0[28] : \regs[11] [28];   // regs.v(45)
    assign n745 = n89 ? wd0[27] : \regs[11] [27];   // regs.v(45)
    assign n746 = n89 ? wd0[26] : \regs[11] [26];   // regs.v(45)
    assign n747 = n89 ? wd0[25] : \regs[11] [25];   // regs.v(45)
    assign n748 = n89 ? wd0[24] : \regs[11] [24];   // regs.v(45)
    assign n749 = n89 ? wd0[23] : \regs[11] [23];   // regs.v(45)
    assign n750 = n89 ? wd0[22] : \regs[11] [22];   // regs.v(45)
    assign n751 = n89 ? wd0[21] : \regs[11] [21];   // regs.v(45)
    assign n752 = n89 ? wd0[20] : \regs[11] [20];   // regs.v(45)
    assign n753 = n89 ? wd0[19] : \regs[11] [19];   // regs.v(45)
    assign n754 = n89 ? wd0[18] : \regs[11] [18];   // regs.v(45)
    assign n755 = n89 ? wd0[17] : \regs[11] [17];   // regs.v(45)
    assign n756 = n89 ? wd0[16] : \regs[11] [16];   // regs.v(45)
    assign n757 = n89 ? wd0[15] : \regs[11] [15];   // regs.v(45)
    assign n758 = n89 ? wd0[14] : \regs[11] [14];   // regs.v(45)
    assign n759 = n89 ? wd0[13] : \regs[11] [13];   // regs.v(45)
    assign n760 = n89 ? wd0[12] : \regs[11] [12];   // regs.v(45)
    assign n761 = n89 ? wd0[11] : \regs[11] [11];   // regs.v(45)
    assign n762 = n89 ? wd0[10] : \regs[11] [10];   // regs.v(45)
    assign n763 = n89 ? wd0[9] : \regs[11] [9];   // regs.v(45)
    assign n764 = n89 ? wd0[8] : \regs[11] [8];   // regs.v(45)
    assign n765 = n89 ? wd0[7] : \regs[11] [7];   // regs.v(45)
    assign n766 = n89 ? wd0[6] : \regs[11] [6];   // regs.v(45)
    assign n767 = n89 ? wd0[5] : \regs[11] [5];   // regs.v(45)
    assign n768 = n89 ? wd0[4] : \regs[11] [4];   // regs.v(45)
    assign n769 = n89 ? wd0[3] : \regs[11] [3];   // regs.v(45)
    assign n770 = n89 ? wd0[2] : \regs[11] [2];   // regs.v(45)
    assign n771 = n89 ? wd0[1] : \regs[11] [1];   // regs.v(45)
    assign n772 = n89 ? wd0[0] : \regs[11] [0];   // regs.v(45)
    assign n773 = n90 ? wd0[31] : \regs[10] [31];   // regs.v(45)
    assign n774 = n90 ? wd0[30] : \regs[10] [30];   // regs.v(45)
    assign n775 = n90 ? wd0[29] : \regs[10] [29];   // regs.v(45)
    assign n776 = n90 ? wd0[28] : \regs[10] [28];   // regs.v(45)
    assign n777 = n90 ? wd0[27] : \regs[10] [27];   // regs.v(45)
    assign n778 = n90 ? wd0[26] : \regs[10] [26];   // regs.v(45)
    assign n779 = n90 ? wd0[25] : \regs[10] [25];   // regs.v(45)
    assign n780 = n90 ? wd0[24] : \regs[10] [24];   // regs.v(45)
    assign n781 = n90 ? wd0[23] : \regs[10] [23];   // regs.v(45)
    assign n782 = n90 ? wd0[22] : \regs[10] [22];   // regs.v(45)
    assign n783 = n90 ? wd0[21] : \regs[10] [21];   // regs.v(45)
    assign n784 = n90 ? wd0[20] : \regs[10] [20];   // regs.v(45)
    assign n785 = n90 ? wd0[19] : \regs[10] [19];   // regs.v(45)
    assign n786 = n90 ? wd0[18] : \regs[10] [18];   // regs.v(45)
    assign n787 = n90 ? wd0[17] : \regs[10] [17];   // regs.v(45)
    assign n788 = n90 ? wd0[16] : \regs[10] [16];   // regs.v(45)
    assign n789 = n90 ? wd0[15] : \regs[10] [15];   // regs.v(45)
    assign n790 = n90 ? wd0[14] : \regs[10] [14];   // regs.v(45)
    assign n791 = n90 ? wd0[13] : \regs[10] [13];   // regs.v(45)
    assign n792 = n90 ? wd0[12] : \regs[10] [12];   // regs.v(45)
    assign n793 = n90 ? wd0[11] : \regs[10] [11];   // regs.v(45)
    assign n794 = n90 ? wd0[10] : \regs[10] [10];   // regs.v(45)
    assign n795 = n90 ? wd0[9] : \regs[10] [9];   // regs.v(45)
    assign n796 = n90 ? wd0[8] : \regs[10] [8];   // regs.v(45)
    assign n797 = n90 ? wd0[7] : \regs[10] [7];   // regs.v(45)
    assign n798 = n90 ? wd0[6] : \regs[10] [6];   // regs.v(45)
    assign n799 = n90 ? wd0[5] : \regs[10] [5];   // regs.v(45)
    assign n800 = n90 ? wd0[4] : \regs[10] [4];   // regs.v(45)
    assign n801 = n90 ? wd0[3] : \regs[10] [3];   // regs.v(45)
    assign n802 = n90 ? wd0[2] : \regs[10] [2];   // regs.v(45)
    assign n803 = n90 ? wd0[1] : \regs[10] [1];   // regs.v(45)
    assign n804 = n90 ? wd0[0] : \regs[10] [0];   // regs.v(45)
    assign n805 = n91 ? wd0[31] : \regs[9] [31];   // regs.v(45)
    assign n806 = n91 ? wd0[30] : \regs[9] [30];   // regs.v(45)
    assign n807 = n91 ? wd0[29] : \regs[9] [29];   // regs.v(45)
    assign n808 = n91 ? wd0[28] : \regs[9] [28];   // regs.v(45)
    assign n809 = n91 ? wd0[27] : \regs[9] [27];   // regs.v(45)
    assign n810 = n91 ? wd0[26] : \regs[9] [26];   // regs.v(45)
    assign n811 = n91 ? wd0[25] : \regs[9] [25];   // regs.v(45)
    assign n812 = n91 ? wd0[24] : \regs[9] [24];   // regs.v(45)
    assign n813 = n91 ? wd0[23] : \regs[9] [23];   // regs.v(45)
    assign n814 = n91 ? wd0[22] : \regs[9] [22];   // regs.v(45)
    assign n815 = n91 ? wd0[21] : \regs[9] [21];   // regs.v(45)
    assign n816 = n91 ? wd0[20] : \regs[9] [20];   // regs.v(45)
    assign n817 = n91 ? wd0[19] : \regs[9] [19];   // regs.v(45)
    assign n818 = n91 ? wd0[18] : \regs[9] [18];   // regs.v(45)
    assign n819 = n91 ? wd0[17] : \regs[9] [17];   // regs.v(45)
    assign n820 = n91 ? wd0[16] : \regs[9] [16];   // regs.v(45)
    assign n821 = n91 ? wd0[15] : \regs[9] [15];   // regs.v(45)
    assign n822 = n91 ? wd0[14] : \regs[9] [14];   // regs.v(45)
    assign n823 = n91 ? wd0[13] : \regs[9] [13];   // regs.v(45)
    assign n824 = n91 ? wd0[12] : \regs[9] [12];   // regs.v(45)
    assign n825 = n91 ? wd0[11] : \regs[9] [11];   // regs.v(45)
    assign n826 = n91 ? wd0[10] : \regs[9] [10];   // regs.v(45)
    assign n827 = n91 ? wd0[9] : \regs[9] [9];   // regs.v(45)
    assign n828 = n91 ? wd0[8] : \regs[9] [8];   // regs.v(45)
    assign n829 = n91 ? wd0[7] : \regs[9] [7];   // regs.v(45)
    assign n830 = n91 ? wd0[6] : \regs[9] [6];   // regs.v(45)
    assign n831 = n91 ? wd0[5] : \regs[9] [5];   // regs.v(45)
    assign n832 = n91 ? wd0[4] : \regs[9] [4];   // regs.v(45)
    assign n833 = n91 ? wd0[3] : \regs[9] [3];   // regs.v(45)
    assign n834 = n91 ? wd0[2] : \regs[9] [2];   // regs.v(45)
    assign n835 = n91 ? wd0[1] : \regs[9] [1];   // regs.v(45)
    assign n836 = n91 ? wd0[0] : \regs[9] [0];   // regs.v(45)
    assign n837 = n92 ? wd0[31] : \regs[8] [31];   // regs.v(45)
    assign n838 = n92 ? wd0[30] : \regs[8] [30];   // regs.v(45)
    assign n839 = n92 ? wd0[29] : \regs[8] [29];   // regs.v(45)
    assign n840 = n92 ? wd0[28] : \regs[8] [28];   // regs.v(45)
    assign n841 = n92 ? wd0[27] : \regs[8] [27];   // regs.v(45)
    assign n842 = n92 ? wd0[26] : \regs[8] [26];   // regs.v(45)
    assign n843 = n92 ? wd0[25] : \regs[8] [25];   // regs.v(45)
    assign n844 = n92 ? wd0[24] : \regs[8] [24];   // regs.v(45)
    assign n845 = n92 ? wd0[23] : \regs[8] [23];   // regs.v(45)
    assign n846 = n92 ? wd0[22] : \regs[8] [22];   // regs.v(45)
    assign n847 = n92 ? wd0[21] : \regs[8] [21];   // regs.v(45)
    assign n848 = n92 ? wd0[20] : \regs[8] [20];   // regs.v(45)
    assign n849 = n92 ? wd0[19] : \regs[8] [19];   // regs.v(45)
    assign n850 = n92 ? wd0[18] : \regs[8] [18];   // regs.v(45)
    assign n851 = n92 ? wd0[17] : \regs[8] [17];   // regs.v(45)
    assign n852 = n92 ? wd0[16] : \regs[8] [16];   // regs.v(45)
    assign n853 = n92 ? wd0[15] : \regs[8] [15];   // regs.v(45)
    assign n854 = n92 ? wd0[14] : \regs[8] [14];   // regs.v(45)
    assign n855 = n92 ? wd0[13] : \regs[8] [13];   // regs.v(45)
    assign n856 = n92 ? wd0[12] : \regs[8] [12];   // regs.v(45)
    assign n857 = n92 ? wd0[11] : \regs[8] [11];   // regs.v(45)
    assign n858 = n92 ? wd0[10] : \regs[8] [10];   // regs.v(45)
    assign n859 = n92 ? wd0[9] : \regs[8] [9];   // regs.v(45)
    assign n860 = n92 ? wd0[8] : \regs[8] [8];   // regs.v(45)
    assign n861 = n92 ? wd0[7] : \regs[8] [7];   // regs.v(45)
    assign n862 = n92 ? wd0[6] : \regs[8] [6];   // regs.v(45)
    assign n863 = n92 ? wd0[5] : \regs[8] [5];   // regs.v(45)
    assign n864 = n92 ? wd0[4] : \regs[8] [4];   // regs.v(45)
    assign n865 = n92 ? wd0[3] : \regs[8] [3];   // regs.v(45)
    assign n866 = n92 ? wd0[2] : \regs[8] [2];   // regs.v(45)
    assign n867 = n92 ? wd0[1] : \regs[8] [1];   // regs.v(45)
    assign n868 = n92 ? wd0[0] : \regs[8] [0];   // regs.v(45)
    assign n869 = n93 ? wd0[31] : \regs[7] [31];   // regs.v(45)
    assign n870 = n93 ? wd0[30] : \regs[7] [30];   // regs.v(45)
    assign n871 = n93 ? wd0[29] : \regs[7] [29];   // regs.v(45)
    assign n872 = n93 ? wd0[28] : \regs[7] [28];   // regs.v(45)
    assign n873 = n93 ? wd0[27] : \regs[7] [27];   // regs.v(45)
    assign n874 = n93 ? wd0[26] : \regs[7] [26];   // regs.v(45)
    assign n875 = n93 ? wd0[25] : \regs[7] [25];   // regs.v(45)
    assign n876 = n93 ? wd0[24] : \regs[7] [24];   // regs.v(45)
    assign n877 = n93 ? wd0[23] : \regs[7] [23];   // regs.v(45)
    assign n878 = n93 ? wd0[22] : \regs[7] [22];   // regs.v(45)
    assign n879 = n93 ? wd0[21] : \regs[7] [21];   // regs.v(45)
    assign n880 = n93 ? wd0[20] : \regs[7] [20];   // regs.v(45)
    assign n881 = n93 ? wd0[19] : \regs[7] [19];   // regs.v(45)
    assign n882 = n93 ? wd0[18] : \regs[7] [18];   // regs.v(45)
    assign n883 = n93 ? wd0[17] : \regs[7] [17];   // regs.v(45)
    assign n884 = n93 ? wd0[16] : \regs[7] [16];   // regs.v(45)
    assign n885 = n93 ? wd0[15] : \regs[7] [15];   // regs.v(45)
    assign n886 = n93 ? wd0[14] : \regs[7] [14];   // regs.v(45)
    assign n887 = n93 ? wd0[13] : \regs[7] [13];   // regs.v(45)
    assign n888 = n93 ? wd0[12] : \regs[7] [12];   // regs.v(45)
    assign n889 = n93 ? wd0[11] : \regs[7] [11];   // regs.v(45)
    assign n890 = n93 ? wd0[10] : \regs[7] [10];   // regs.v(45)
    assign n891 = n93 ? wd0[9] : \regs[7] [9];   // regs.v(45)
    assign n892 = n93 ? wd0[8] : \regs[7] [8];   // regs.v(45)
    assign n893 = n93 ? wd0[7] : \regs[7] [7];   // regs.v(45)
    assign n894 = n93 ? wd0[6] : \regs[7] [6];   // regs.v(45)
    assign n895 = n93 ? wd0[5] : \regs[7] [5];   // regs.v(45)
    assign n896 = n93 ? wd0[4] : \regs[7] [4];   // regs.v(45)
    assign n897 = n93 ? wd0[3] : \regs[7] [3];   // regs.v(45)
    assign n898 = n93 ? wd0[2] : \regs[7] [2];   // regs.v(45)
    assign n899 = n93 ? wd0[1] : \regs[7] [1];   // regs.v(45)
    assign n900 = n93 ? wd0[0] : \regs[7] [0];   // regs.v(45)
    assign n901 = n94 ? wd0[31] : \regs[6] [31];   // regs.v(45)
    assign n902 = n94 ? wd0[30] : \regs[6] [30];   // regs.v(45)
    assign n903 = n94 ? wd0[29] : \regs[6] [29];   // regs.v(45)
    assign n904 = n94 ? wd0[28] : \regs[6] [28];   // regs.v(45)
    assign n905 = n94 ? wd0[27] : \regs[6] [27];   // regs.v(45)
    assign n906 = n94 ? wd0[26] : \regs[6] [26];   // regs.v(45)
    assign n907 = n94 ? wd0[25] : \regs[6] [25];   // regs.v(45)
    assign n908 = n94 ? wd0[24] : \regs[6] [24];   // regs.v(45)
    assign n909 = n94 ? wd0[23] : \regs[6] [23];   // regs.v(45)
    assign n910 = n94 ? wd0[22] : \regs[6] [22];   // regs.v(45)
    assign n911 = n94 ? wd0[21] : \regs[6] [21];   // regs.v(45)
    assign n912 = n94 ? wd0[20] : \regs[6] [20];   // regs.v(45)
    assign n913 = n94 ? wd0[19] : \regs[6] [19];   // regs.v(45)
    assign n914 = n94 ? wd0[18] : \regs[6] [18];   // regs.v(45)
    assign n915 = n94 ? wd0[17] : \regs[6] [17];   // regs.v(45)
    assign n916 = n94 ? wd0[16] : \regs[6] [16];   // regs.v(45)
    assign n917 = n94 ? wd0[15] : \regs[6] [15];   // regs.v(45)
    assign n918 = n94 ? wd0[14] : \regs[6] [14];   // regs.v(45)
    assign n919 = n94 ? wd0[13] : \regs[6] [13];   // regs.v(45)
    assign n920 = n94 ? wd0[12] : \regs[6] [12];   // regs.v(45)
    assign n921 = n94 ? wd0[11] : \regs[6] [11];   // regs.v(45)
    assign n922 = n94 ? wd0[10] : \regs[6] [10];   // regs.v(45)
    assign n923 = n94 ? wd0[9] : \regs[6] [9];   // regs.v(45)
    assign n924 = n94 ? wd0[8] : \regs[6] [8];   // regs.v(45)
    assign n925 = n94 ? wd0[7] : \regs[6] [7];   // regs.v(45)
    assign n926 = n94 ? wd0[6] : \regs[6] [6];   // regs.v(45)
    assign n927 = n94 ? wd0[5] : \regs[6] [5];   // regs.v(45)
    assign n928 = n94 ? wd0[4] : \regs[6] [4];   // regs.v(45)
    assign n929 = n94 ? wd0[3] : \regs[6] [3];   // regs.v(45)
    assign n930 = n94 ? wd0[2] : \regs[6] [2];   // regs.v(45)
    assign n931 = n94 ? wd0[1] : \regs[6] [1];   // regs.v(45)
    assign n932 = n94 ? wd0[0] : \regs[6] [0];   // regs.v(45)
    assign n933 = n95 ? wd0[31] : \regs[5] [31];   // regs.v(45)
    assign n934 = n95 ? wd0[30] : \regs[5] [30];   // regs.v(45)
    assign n935 = n95 ? wd0[29] : \regs[5] [29];   // regs.v(45)
    assign n936 = n95 ? wd0[28] : \regs[5] [28];   // regs.v(45)
    assign n937 = n95 ? wd0[27] : \regs[5] [27];   // regs.v(45)
    assign n938 = n95 ? wd0[26] : \regs[5] [26];   // regs.v(45)
    assign n939 = n95 ? wd0[25] : \regs[5] [25];   // regs.v(45)
    assign n940 = n95 ? wd0[24] : \regs[5] [24];   // regs.v(45)
    assign n941 = n95 ? wd0[23] : \regs[5] [23];   // regs.v(45)
    assign n942 = n95 ? wd0[22] : \regs[5] [22];   // regs.v(45)
    assign n943 = n95 ? wd0[21] : \regs[5] [21];   // regs.v(45)
    assign n944 = n95 ? wd0[20] : \regs[5] [20];   // regs.v(45)
    assign n945 = n95 ? wd0[19] : \regs[5] [19];   // regs.v(45)
    assign n946 = n95 ? wd0[18] : \regs[5] [18];   // regs.v(45)
    assign n947 = n95 ? wd0[17] : \regs[5] [17];   // regs.v(45)
    assign n948 = n95 ? wd0[16] : \regs[5] [16];   // regs.v(45)
    assign n949 = n95 ? wd0[15] : \regs[5] [15];   // regs.v(45)
    assign n950 = n95 ? wd0[14] : \regs[5] [14];   // regs.v(45)
    assign n951 = n95 ? wd0[13] : \regs[5] [13];   // regs.v(45)
    assign n952 = n95 ? wd0[12] : \regs[5] [12];   // regs.v(45)
    assign n953 = n95 ? wd0[11] : \regs[5] [11];   // regs.v(45)
    assign n954 = n95 ? wd0[10] : \regs[5] [10];   // regs.v(45)
    assign n955 = n95 ? wd0[9] : \regs[5] [9];   // regs.v(45)
    assign n956 = n95 ? wd0[8] : \regs[5] [8];   // regs.v(45)
    assign n957 = n95 ? wd0[7] : \regs[5] [7];   // regs.v(45)
    assign n958 = n95 ? wd0[6] : \regs[5] [6];   // regs.v(45)
    assign n959 = n95 ? wd0[5] : \regs[5] [5];   // regs.v(45)
    assign n960 = n95 ? wd0[4] : \regs[5] [4];   // regs.v(45)
    assign n961 = n95 ? wd0[3] : \regs[5] [3];   // regs.v(45)
    assign n962 = n95 ? wd0[2] : \regs[5] [2];   // regs.v(45)
    assign n963 = n95 ? wd0[1] : \regs[5] [1];   // regs.v(45)
    assign n964 = n95 ? wd0[0] : \regs[5] [0];   // regs.v(45)
    assign n965 = n96 ? wd0[31] : \regs[4] [31];   // regs.v(45)
    assign n966 = n96 ? wd0[30] : \regs[4] [30];   // regs.v(45)
    assign n967 = n96 ? wd0[29] : \regs[4] [29];   // regs.v(45)
    assign n968 = n96 ? wd0[28] : \regs[4] [28];   // regs.v(45)
    assign n969 = n96 ? wd0[27] : \regs[4] [27];   // regs.v(45)
    assign n970 = n96 ? wd0[26] : \regs[4] [26];   // regs.v(45)
    assign n971 = n96 ? wd0[25] : \regs[4] [25];   // regs.v(45)
    assign n972 = n96 ? wd0[24] : \regs[4] [24];   // regs.v(45)
    assign n973 = n96 ? wd0[23] : \regs[4] [23];   // regs.v(45)
    assign n974 = n96 ? wd0[22] : \regs[4] [22];   // regs.v(45)
    assign n975 = n96 ? wd0[21] : \regs[4] [21];   // regs.v(45)
    assign n976 = n96 ? wd0[20] : \regs[4] [20];   // regs.v(45)
    assign n977 = n96 ? wd0[19] : \regs[4] [19];   // regs.v(45)
    assign n978 = n96 ? wd0[18] : \regs[4] [18];   // regs.v(45)
    assign n979 = n96 ? wd0[17] : \regs[4] [17];   // regs.v(45)
    assign n980 = n96 ? wd0[16] : \regs[4] [16];   // regs.v(45)
    assign n981 = n96 ? wd0[15] : \regs[4] [15];   // regs.v(45)
    assign n982 = n96 ? wd0[14] : \regs[4] [14];   // regs.v(45)
    assign n983 = n96 ? wd0[13] : \regs[4] [13];   // regs.v(45)
    assign n984 = n96 ? wd0[12] : \regs[4] [12];   // regs.v(45)
    assign n985 = n96 ? wd0[11] : \regs[4] [11];   // regs.v(45)
    assign n986 = n96 ? wd0[10] : \regs[4] [10];   // regs.v(45)
    assign n987 = n96 ? wd0[9] : \regs[4] [9];   // regs.v(45)
    assign n988 = n96 ? wd0[8] : \regs[4] [8];   // regs.v(45)
    assign n989 = n96 ? wd0[7] : \regs[4] [7];   // regs.v(45)
    assign n990 = n96 ? wd0[6] : \regs[4] [6];   // regs.v(45)
    assign n991 = n96 ? wd0[5] : \regs[4] [5];   // regs.v(45)
    assign n992 = n96 ? wd0[4] : \regs[4] [4];   // regs.v(45)
    assign n993 = n96 ? wd0[3] : \regs[4] [3];   // regs.v(45)
    assign n994 = n96 ? wd0[2] : \regs[4] [2];   // regs.v(45)
    assign n995 = n96 ? wd0[1] : \regs[4] [1];   // regs.v(45)
    assign n996 = n96 ? wd0[0] : \regs[4] [0];   // regs.v(45)
    assign n997 = n97 ? wd0[31] : \regs[3] [31];   // regs.v(45)
    assign n998 = n97 ? wd0[30] : \regs[3] [30];   // regs.v(45)
    assign n999 = n97 ? wd0[29] : \regs[3] [29];   // regs.v(45)
    assign n1000 = n97 ? wd0[28] : \regs[3] [28];   // regs.v(45)
    assign n1001 = n97 ? wd0[27] : \regs[3] [27];   // regs.v(45)
    assign n1002 = n97 ? wd0[26] : \regs[3] [26];   // regs.v(45)
    assign n1003 = n97 ? wd0[25] : \regs[3] [25];   // regs.v(45)
    assign n1004 = n97 ? wd0[24] : \regs[3] [24];   // regs.v(45)
    assign n1005 = n97 ? wd0[23] : \regs[3] [23];   // regs.v(45)
    assign n1006 = n97 ? wd0[22] : \regs[3] [22];   // regs.v(45)
    assign n1007 = n97 ? wd0[21] : \regs[3] [21];   // regs.v(45)
    assign n1008 = n97 ? wd0[20] : \regs[3] [20];   // regs.v(45)
    assign n1009 = n97 ? wd0[19] : \regs[3] [19];   // regs.v(45)
    assign n1010 = n97 ? wd0[18] : \regs[3] [18];   // regs.v(45)
    assign n1011 = n97 ? wd0[17] : \regs[3] [17];   // regs.v(45)
    assign n1012 = n97 ? wd0[16] : \regs[3] [16];   // regs.v(45)
    assign n1013 = n97 ? wd0[15] : \regs[3] [15];   // regs.v(45)
    assign n1014 = n97 ? wd0[14] : \regs[3] [14];   // regs.v(45)
    assign n1015 = n97 ? wd0[13] : \regs[3] [13];   // regs.v(45)
    assign n1016 = n97 ? wd0[12] : \regs[3] [12];   // regs.v(45)
    assign n1017 = n97 ? wd0[11] : \regs[3] [11];   // regs.v(45)
    assign n1018 = n97 ? wd0[10] : \regs[3] [10];   // regs.v(45)
    assign n1019 = n97 ? wd0[9] : \regs[3] [9];   // regs.v(45)
    assign n1020 = n97 ? wd0[8] : \regs[3] [8];   // regs.v(45)
    assign n1021 = n97 ? wd0[7] : \regs[3] [7];   // regs.v(45)
    assign n1022 = n97 ? wd0[6] : \regs[3] [6];   // regs.v(45)
    assign n1023 = n97 ? wd0[5] : \regs[3] [5];   // regs.v(45)
    assign n1024 = n97 ? wd0[4] : \regs[3] [4];   // regs.v(45)
    assign n1025 = n97 ? wd0[3] : \regs[3] [3];   // regs.v(45)
    assign n1026 = n97 ? wd0[2] : \regs[3] [2];   // regs.v(45)
    assign n1027 = n97 ? wd0[1] : \regs[3] [1];   // regs.v(45)
    assign n1028 = n97 ? wd0[0] : \regs[3] [0];   // regs.v(45)
    assign n1029 = n98 ? wd0[31] : \regs[2] [31];   // regs.v(45)
    assign n1030 = n98 ? wd0[30] : \regs[2] [30];   // regs.v(45)
    assign n1031 = n98 ? wd0[29] : \regs[2] [29];   // regs.v(45)
    assign n1032 = n98 ? wd0[28] : \regs[2] [28];   // regs.v(45)
    assign n1033 = n98 ? wd0[27] : \regs[2] [27];   // regs.v(45)
    assign n1034 = n98 ? wd0[26] : \regs[2] [26];   // regs.v(45)
    assign n1035 = n98 ? wd0[25] : \regs[2] [25];   // regs.v(45)
    assign n1036 = n98 ? wd0[24] : \regs[2] [24];   // regs.v(45)
    assign n1037 = n98 ? wd0[23] : \regs[2] [23];   // regs.v(45)
    assign n1038 = n98 ? wd0[22] : \regs[2] [22];   // regs.v(45)
    assign n1039 = n98 ? wd0[21] : \regs[2] [21];   // regs.v(45)
    assign n1040 = n98 ? wd0[20] : \regs[2] [20];   // regs.v(45)
    assign n1041 = n98 ? wd0[19] : \regs[2] [19];   // regs.v(45)
    assign n1042 = n98 ? wd0[18] : \regs[2] [18];   // regs.v(45)
    assign n1043 = n98 ? wd0[17] : \regs[2] [17];   // regs.v(45)
    assign n1044 = n98 ? wd0[16] : \regs[2] [16];   // regs.v(45)
    assign n1045 = n98 ? wd0[15] : \regs[2] [15];   // regs.v(45)
    assign n1046 = n98 ? wd0[14] : \regs[2] [14];   // regs.v(45)
    assign n1047 = n98 ? wd0[13] : \regs[2] [13];   // regs.v(45)
    assign n1048 = n98 ? wd0[12] : \regs[2] [12];   // regs.v(45)
    assign n1049 = n98 ? wd0[11] : \regs[2] [11];   // regs.v(45)
    assign n1050 = n98 ? wd0[10] : \regs[2] [10];   // regs.v(45)
    assign n1051 = n98 ? wd0[9] : \regs[2] [9];   // regs.v(45)
    assign n1052 = n98 ? wd0[8] : \regs[2] [8];   // regs.v(45)
    assign n1053 = n98 ? wd0[7] : \regs[2] [7];   // regs.v(45)
    assign n1054 = n98 ? wd0[6] : \regs[2] [6];   // regs.v(45)
    assign n1055 = n98 ? wd0[5] : \regs[2] [5];   // regs.v(45)
    assign n1056 = n98 ? wd0[4] : \regs[2] [4];   // regs.v(45)
    assign n1057 = n98 ? wd0[3] : \regs[2] [3];   // regs.v(45)
    assign n1058 = n98 ? wd0[2] : \regs[2] [2];   // regs.v(45)
    assign n1059 = n98 ? wd0[1] : \regs[2] [1];   // regs.v(45)
    assign n1060 = n98 ? wd0[0] : \regs[2] [0];   // regs.v(45)
    assign n1061 = n99 ? wd0[31] : \regs[1] [31];   // regs.v(45)
    assign n1062 = n99 ? wd0[30] : \regs[1] [30];   // regs.v(45)
    assign n1063 = n99 ? wd0[29] : \regs[1] [29];   // regs.v(45)
    assign n1064 = n99 ? wd0[28] : \regs[1] [28];   // regs.v(45)
    assign n1065 = n99 ? wd0[27] : \regs[1] [27];   // regs.v(45)
    assign n1066 = n99 ? wd0[26] : \regs[1] [26];   // regs.v(45)
    assign n1067 = n99 ? wd0[25] : \regs[1] [25];   // regs.v(45)
    assign n1068 = n99 ? wd0[24] : \regs[1] [24];   // regs.v(45)
    assign n1069 = n99 ? wd0[23] : \regs[1] [23];   // regs.v(45)
    assign n1070 = n99 ? wd0[22] : \regs[1] [22];   // regs.v(45)
    assign n1071 = n99 ? wd0[21] : \regs[1] [21];   // regs.v(45)
    assign n1072 = n99 ? wd0[20] : \regs[1] [20];   // regs.v(45)
    assign n1073 = n99 ? wd0[19] : \regs[1] [19];   // regs.v(45)
    assign n1074 = n99 ? wd0[18] : \regs[1] [18];   // regs.v(45)
    assign n1075 = n99 ? wd0[17] : \regs[1] [17];   // regs.v(45)
    assign n1076 = n99 ? wd0[16] : \regs[1] [16];   // regs.v(45)
    assign n1077 = n99 ? wd0[15] : \regs[1] [15];   // regs.v(45)
    assign n1078 = n99 ? wd0[14] : \regs[1] [14];   // regs.v(45)
    assign n1079 = n99 ? wd0[13] : \regs[1] [13];   // regs.v(45)
    assign n1080 = n99 ? wd0[12] : \regs[1] [12];   // regs.v(45)
    assign n1081 = n99 ? wd0[11] : \regs[1] [11];   // regs.v(45)
    assign n1082 = n99 ? wd0[10] : \regs[1] [10];   // regs.v(45)
    assign n1083 = n99 ? wd0[9] : \regs[1] [9];   // regs.v(45)
    assign n1084 = n99 ? wd0[8] : \regs[1] [8];   // regs.v(45)
    assign n1085 = n99 ? wd0[7] : \regs[1] [7];   // regs.v(45)
    assign n1086 = n99 ? wd0[6] : \regs[1] [6];   // regs.v(45)
    assign n1087 = n99 ? wd0[5] : \regs[1] [5];   // regs.v(45)
    assign n1088 = n99 ? wd0[4] : \regs[1] [4];   // regs.v(45)
    assign n1089 = n99 ? wd0[3] : \regs[1] [3];   // regs.v(45)
    assign n1090 = n99 ? wd0[2] : \regs[1] [2];   // regs.v(45)
    assign n1091 = n99 ? wd0[1] : \regs[1] [1];   // regs.v(45)
    assign n1092 = n99 ? wd0[0] : \regs[1] [0];   // regs.v(45)
    assign n1093 = n100 ? wd0[31] : \regs[0] [31];   // regs.v(45)
    assign n1094 = n100 ? wd0[30] : \regs[0] [30];   // regs.v(45)
    assign n1095 = n100 ? wd0[29] : \regs[0] [29];   // regs.v(45)
    assign n1096 = n100 ? wd0[28] : \regs[0] [28];   // regs.v(45)
    assign n1097 = n100 ? wd0[27] : \regs[0] [27];   // regs.v(45)
    assign n1098 = n100 ? wd0[26] : \regs[0] [26];   // regs.v(45)
    assign n1099 = n100 ? wd0[25] : \regs[0] [25];   // regs.v(45)
    assign n1100 = n100 ? wd0[24] : \regs[0] [24];   // regs.v(45)
    assign n1101 = n100 ? wd0[23] : \regs[0] [23];   // regs.v(45)
    assign n1102 = n100 ? wd0[22] : \regs[0] [22];   // regs.v(45)
    assign n1103 = n100 ? wd0[21] : \regs[0] [21];   // regs.v(45)
    assign n1104 = n100 ? wd0[20] : \regs[0] [20];   // regs.v(45)
    assign n1105 = n100 ? wd0[19] : \regs[0] [19];   // regs.v(45)
    assign n1106 = n100 ? wd0[18] : \regs[0] [18];   // regs.v(45)
    assign n1107 = n100 ? wd0[17] : \regs[0] [17];   // regs.v(45)
    assign n1108 = n100 ? wd0[16] : \regs[0] [16];   // regs.v(45)
    assign n1109 = n100 ? wd0[15] : \regs[0] [15];   // regs.v(45)
    assign n1110 = n100 ? wd0[14] : \regs[0] [14];   // regs.v(45)
    assign n1111 = n100 ? wd0[13] : \regs[0] [13];   // regs.v(45)
    assign n1112 = n100 ? wd0[12] : \regs[0] [12];   // regs.v(45)
    assign n1113 = n100 ? wd0[11] : \regs[0] [11];   // regs.v(45)
    assign n1114 = n100 ? wd0[10] : \regs[0] [10];   // regs.v(45)
    assign n1115 = n100 ? wd0[9] : \regs[0] [9];   // regs.v(45)
    assign n1116 = n100 ? wd0[8] : \regs[0] [8];   // regs.v(45)
    assign n1117 = n100 ? wd0[7] : \regs[0] [7];   // regs.v(45)
    assign n1118 = n100 ? wd0[6] : \regs[0] [6];   // regs.v(45)
    assign n1119 = n100 ? wd0[5] : \regs[0] [5];   // regs.v(45)
    assign n1120 = n100 ? wd0[4] : \regs[0] [4];   // regs.v(45)
    assign n1121 = n100 ? wd0[3] : \regs[0] [3];   // regs.v(45)
    assign n1122 = n100 ? wd0[2] : \regs[0] [2];   // regs.v(45)
    assign n1123 = n100 ? wd0[1] : \regs[0] [1];   // regs.v(45)
    assign n1124 = n100 ? wd0[0] : \regs[0] [0];   // regs.v(45)
    assign n1125 = write[0] ? n101 : pcout[31];   // regs.v(45)
    assign n1126 = write[0] ? n102 : pcout[30];   // regs.v(45)
    assign n1127 = write[0] ? n103 : pcout[29];   // regs.v(45)
    assign n1128 = write[0] ? n104 : pcout[28];   // regs.v(45)
    assign n1129 = write[0] ? n105 : pcout[27];   // regs.v(45)
    assign n1130 = write[0] ? n106 : pcout[26];   // regs.v(45)
    assign n1131 = write[0] ? n107 : pcout[25];   // regs.v(45)
    assign n1132 = write[0] ? n108 : pcout[24];   // regs.v(45)
    assign n1133 = write[0] ? n109 : pcout[23];   // regs.v(45)
    assign n1134 = write[0] ? n110 : pcout[22];   // regs.v(45)
    assign n1135 = write[0] ? n111 : pcout[21];   // regs.v(45)
    assign n1136 = write[0] ? n112 : pcout[20];   // regs.v(45)
    assign n1137 = write[0] ? n113 : pcout[19];   // regs.v(45)
    assign n1138 = write[0] ? n114 : pcout[18];   // regs.v(45)
    assign n1139 = write[0] ? n115 : pcout[17];   // regs.v(45)
    assign n1140 = write[0] ? n116 : pcout[16];   // regs.v(45)
    assign n1141 = write[0] ? n117 : pcout[15];   // regs.v(45)
    assign n1142 = write[0] ? n118 : pcout[14];   // regs.v(45)
    assign n1143 = write[0] ? n119 : pcout[13];   // regs.v(45)
    assign n1144 = write[0] ? n120 : pcout[12];   // regs.v(45)
    assign n1145 = write[0] ? n121 : pcout[11];   // regs.v(45)
    assign n1146 = write[0] ? n122 : pcout[10];   // regs.v(45)
    assign n1147 = write[0] ? n123 : pcout[9];   // regs.v(45)
    assign n1148 = write[0] ? n124 : pcout[8];   // regs.v(45)
    assign n1149 = write[0] ? n125 : pcout[7];   // regs.v(45)
    assign n1150 = write[0] ? n126 : pcout[6];   // regs.v(45)
    assign n1151 = write[0] ? n127 : pcout[5];   // regs.v(45)
    assign n1152 = write[0] ? n128 : pcout[4];   // regs.v(45)
    assign n1153 = write[0] ? n129 : pcout[3];   // regs.v(45)
    assign n1154 = write[0] ? n130 : pcout[2];   // regs.v(45)
    assign n1155 = write[0] ? n131 : pcout[1];   // regs.v(45)
    assign n1156 = write[0] ? n132 : pcout[0];   // regs.v(45)
    assign n1157 = write[0] ? n133 : spout[31];   // regs.v(45)
    assign n1158 = write[0] ? n134 : spout[30];   // regs.v(45)
    assign n1159 = write[0] ? n135 : spout[29];   // regs.v(45)
    assign n1160 = write[0] ? n136 : spout[28];   // regs.v(45)
    assign n1161 = write[0] ? n137 : spout[27];   // regs.v(45)
    assign n1162 = write[0] ? n138 : spout[26];   // regs.v(45)
    assign n1163 = write[0] ? n139 : spout[25];   // regs.v(45)
    assign n1164 = write[0] ? n140 : spout[24];   // regs.v(45)
    assign n1165 = write[0] ? n141 : spout[23];   // regs.v(45)
    assign n1166 = write[0] ? n142 : spout[22];   // regs.v(45)
    assign n1167 = write[0] ? n143 : spout[21];   // regs.v(45)
    assign n1168 = write[0] ? n144 : spout[20];   // regs.v(45)
    assign n1169 = write[0] ? n145 : spout[19];   // regs.v(45)
    assign n1170 = write[0] ? n146 : spout[18];   // regs.v(45)
    assign n1171 = write[0] ? n147 : spout[17];   // regs.v(45)
    assign n1172 = write[0] ? n148 : spout[16];   // regs.v(45)
    assign n1173 = write[0] ? n149 : spout[15];   // regs.v(45)
    assign n1174 = write[0] ? n150 : spout[14];   // regs.v(45)
    assign n1175 = write[0] ? n151 : spout[13];   // regs.v(45)
    assign n1176 = write[0] ? n152 : spout[12];   // regs.v(45)
    assign n1177 = write[0] ? n153 : spout[11];   // regs.v(45)
    assign n1178 = write[0] ? n154 : spout[10];   // regs.v(45)
    assign n1179 = write[0] ? n155 : spout[9];   // regs.v(45)
    assign n1180 = write[0] ? n156 : spout[8];   // regs.v(45)
    assign n1181 = write[0] ? n157 : spout[7];   // regs.v(45)
    assign n1182 = write[0] ? n158 : spout[6];   // regs.v(45)
    assign n1183 = write[0] ? n159 : spout[5];   // regs.v(45)
    assign n1184 = write[0] ? n160 : spout[4];   // regs.v(45)
    assign n1185 = write[0] ? n161 : spout[3];   // regs.v(45)
    assign n1186 = write[0] ? n162 : spout[2];   // regs.v(45)
    assign n1187 = write[0] ? n163 : spout[1];   // regs.v(45)
    assign n1188 = write[0] ? n164 : spout[0];   // regs.v(45)
    assign n1189 = write[0] ? n165 : lrout[31];   // regs.v(45)
    assign n1190 = write[0] ? n166 : lrout[30];   // regs.v(45)
    assign n1191 = write[0] ? n167 : lrout[29];   // regs.v(45)
    assign n1192 = write[0] ? n168 : lrout[28];   // regs.v(45)
    assign n1193 = write[0] ? n169 : lrout[27];   // regs.v(45)
    assign n1194 = write[0] ? n170 : lrout[26];   // regs.v(45)
    assign n1195 = write[0] ? n171 : lrout[25];   // regs.v(45)
    assign n1196 = write[0] ? n172 : lrout[24];   // regs.v(45)
    assign n1197 = write[0] ? n173 : lrout[23];   // regs.v(45)
    assign n1198 = write[0] ? n174 : lrout[22];   // regs.v(45)
    assign n1199 = write[0] ? n175 : lrout[21];   // regs.v(45)
    assign n1200 = write[0] ? n176 : lrout[20];   // regs.v(45)
    assign n1201 = write[0] ? n177 : lrout[19];   // regs.v(45)
    assign n1202 = write[0] ? n178 : lrout[18];   // regs.v(45)
    assign n1203 = write[0] ? n179 : lrout[17];   // regs.v(45)
    assign n1204 = write[0] ? n180 : lrout[16];   // regs.v(45)
    assign n1205 = write[0] ? n181 : lrout[15];   // regs.v(45)
    assign n1206 = write[0] ? n182 : lrout[14];   // regs.v(45)
    assign n1207 = write[0] ? n183 : lrout[13];   // regs.v(45)
    assign n1208 = write[0] ? n184 : lrout[12];   // regs.v(45)
    assign n1209 = write[0] ? n185 : lrout[11];   // regs.v(45)
    assign n1210 = write[0] ? n186 : lrout[10];   // regs.v(45)
    assign n1211 = write[0] ? n187 : lrout[9];   // regs.v(45)
    assign n1212 = write[0] ? n188 : lrout[8];   // regs.v(45)
    assign n1213 = write[0] ? n189 : lrout[7];   // regs.v(45)
    assign n1214 = write[0] ? n190 : lrout[6];   // regs.v(45)
    assign n1215 = write[0] ? n191 : lrout[5];   // regs.v(45)
    assign n1216 = write[0] ? n192 : lrout[4];   // regs.v(45)
    assign n1217 = write[0] ? n193 : lrout[3];   // regs.v(45)
    assign n1218 = write[0] ? n194 : lrout[2];   // regs.v(45)
    assign n1219 = write[0] ? n195 : lrout[1];   // regs.v(45)
    assign n1220 = write[0] ? n196 : lrout[0];   // regs.v(45)
    assign n1221 = write[0] ? n197 : stout[31];   // regs.v(45)
    assign n1222 = write[0] ? n198 : stout[30];   // regs.v(45)
    assign n1223 = write[0] ? n199 : stout[29];   // regs.v(45)
    assign n1224 = write[0] ? n200 : stout[28];   // regs.v(45)
    assign n1225 = write[0] ? n201 : stout[27];   // regs.v(45)
    assign n1226 = write[0] ? n202 : stout[26];   // regs.v(45)
    assign n1227 = write[0] ? n203 : stout[25];   // regs.v(45)
    assign n1228 = write[0] ? n204 : stout[24];   // regs.v(45)
    assign n1229 = write[0] ? n205 : stout[23];   // regs.v(45)
    assign n1230 = write[0] ? n206 : stout[22];   // regs.v(45)
    assign n1231 = write[0] ? n207 : stout[21];   // regs.v(45)
    assign n1232 = write[0] ? n208 : stout[20];   // regs.v(45)
    assign n1233 = write[0] ? n209 : stout[19];   // regs.v(45)
    assign n1234 = write[0] ? n210 : stout[18];   // regs.v(45)
    assign n1235 = write[0] ? n211 : stout[17];   // regs.v(45)
    assign n1236 = write[0] ? n212 : stout[16];   // regs.v(45)
    assign n1237 = write[0] ? n213 : stout[15];   // regs.v(45)
    assign n1238 = write[0] ? n214 : stout[14];   // regs.v(45)
    assign n1239 = write[0] ? n215 : stout[13];   // regs.v(45)
    assign n1240 = write[0] ? n216 : stout[12];   // regs.v(45)
    assign n1241 = write[0] ? n217 : stout[11];   // regs.v(45)
    assign n1242 = write[0] ? n218 : stout[10];   // regs.v(45)
    assign n1243 = write[0] ? n219 : stout[9];   // regs.v(45)
    assign n1244 = write[0] ? n220 : stout[8];   // regs.v(45)
    assign n1245 = write[0] ? n221 : stout[7];   // regs.v(45)
    assign n1246 = write[0] ? n222 : stout[6];   // regs.v(45)
    assign n1247 = write[0] ? n223 : stout[5];   // regs.v(45)
    assign n1248 = write[0] ? n224 : stout[4];   // regs.v(45)
    assign n1249 = write[0] ? n225 : stout[3];   // regs.v(45)
    assign n1250 = write[0] ? n226 : stout[2];   // regs.v(45)
    assign n1251 = write[0] ? n227 : stout[1];   // regs.v(45)
    assign n1252 = write[0] ? n228 : stout[0];   // regs.v(45)
    assign n1253 = write[0] ? n229 : \regs[27] [31];   // regs.v(45)
    assign n1254 = write[0] ? n230 : \regs[27] [30];   // regs.v(45)
    assign n1255 = write[0] ? n231 : \regs[27] [29];   // regs.v(45)
    assign n1256 = write[0] ? n232 : \regs[27] [28];   // regs.v(45)
    assign n1257 = write[0] ? n233 : \regs[27] [27];   // regs.v(45)
    assign n1258 = write[0] ? n234 : \regs[27] [26];   // regs.v(45)
    assign n1259 = write[0] ? n235 : \regs[27] [25];   // regs.v(45)
    assign n1260 = write[0] ? n236 : \regs[27] [24];   // regs.v(45)
    assign n1261 = write[0] ? n237 : \regs[27] [23];   // regs.v(45)
    assign n1262 = write[0] ? n238 : \regs[27] [22];   // regs.v(45)
    assign n1263 = write[0] ? n239 : \regs[27] [21];   // regs.v(45)
    assign n1264 = write[0] ? n240 : \regs[27] [20];   // regs.v(45)
    assign n1265 = write[0] ? n241 : \regs[27] [19];   // regs.v(45)
    assign n1266 = write[0] ? n242 : \regs[27] [18];   // regs.v(45)
    assign n1267 = write[0] ? n243 : \regs[27] [17];   // regs.v(45)
    assign n1268 = write[0] ? n244 : \regs[27] [16];   // regs.v(45)
    assign n1269 = write[0] ? n245 : \regs[27] [15];   // regs.v(45)
    assign n1270 = write[0] ? n246 : \regs[27] [14];   // regs.v(45)
    assign n1271 = write[0] ? n247 : \regs[27] [13];   // regs.v(45)
    assign n1272 = write[0] ? n248 : \regs[27] [12];   // regs.v(45)
    assign n1273 = write[0] ? n249 : \regs[27] [11];   // regs.v(45)
    assign n1274 = write[0] ? n250 : \regs[27] [10];   // regs.v(45)
    assign n1275 = write[0] ? n251 : \regs[27] [9];   // regs.v(45)
    assign n1276 = write[0] ? n252 : \regs[27] [8];   // regs.v(45)
    assign n1277 = write[0] ? n253 : \regs[27] [7];   // regs.v(45)
    assign n1278 = write[0] ? n254 : \regs[27] [6];   // regs.v(45)
    assign n1279 = write[0] ? n255 : \regs[27] [5];   // regs.v(45)
    assign n1280 = write[0] ? n256 : \regs[27] [4];   // regs.v(45)
    assign n1281 = write[0] ? n257 : \regs[27] [3];   // regs.v(45)
    assign n1282 = write[0] ? n258 : \regs[27] [2];   // regs.v(45)
    assign n1283 = write[0] ? n259 : \regs[27] [1];   // regs.v(45)
    assign n1284 = write[0] ? n260 : \regs[27] [0];   // regs.v(45)
    assign n1285 = write[0] ? n261 : \regs[26] [31];   // regs.v(45)
    assign n1286 = write[0] ? n262 : \regs[26] [30];   // regs.v(45)
    assign n1287 = write[0] ? n263 : \regs[26] [29];   // regs.v(45)
    assign n1288 = write[0] ? n264 : \regs[26] [28];   // regs.v(45)
    assign n1289 = write[0] ? n265 : \regs[26] [27];   // regs.v(45)
    assign n1290 = write[0] ? n266 : \regs[26] [26];   // regs.v(45)
    assign n1291 = write[0] ? n267 : \regs[26] [25];   // regs.v(45)
    assign n1292 = write[0] ? n268 : \regs[26] [24];   // regs.v(45)
    assign n1293 = write[0] ? n269 : \regs[26] [23];   // regs.v(45)
    assign n1294 = write[0] ? n270 : \regs[26] [22];   // regs.v(45)
    assign n1295 = write[0] ? n271 : \regs[26] [21];   // regs.v(45)
    assign n1296 = write[0] ? n272 : \regs[26] [20];   // regs.v(45)
    assign n1297 = write[0] ? n273 : \regs[26] [19];   // regs.v(45)
    assign n1298 = write[0] ? n274 : \regs[26] [18];   // regs.v(45)
    assign n1299 = write[0] ? n275 : \regs[26] [17];   // regs.v(45)
    assign n1300 = write[0] ? n276 : \regs[26] [16];   // regs.v(45)
    assign n1301 = write[0] ? n277 : \regs[26] [15];   // regs.v(45)
    assign n1302 = write[0] ? n278 : \regs[26] [14];   // regs.v(45)
    assign n1303 = write[0] ? n279 : \regs[26] [13];   // regs.v(45)
    assign n1304 = write[0] ? n280 : \regs[26] [12];   // regs.v(45)
    assign n1305 = write[0] ? n281 : \regs[26] [11];   // regs.v(45)
    assign n1306 = write[0] ? n282 : \regs[26] [10];   // regs.v(45)
    assign n1307 = write[0] ? n283 : \regs[26] [9];   // regs.v(45)
    assign n1308 = write[0] ? n284 : \regs[26] [8];   // regs.v(45)
    assign n1309 = write[0] ? n285 : \regs[26] [7];   // regs.v(45)
    assign n1310 = write[0] ? n286 : \regs[26] [6];   // regs.v(45)
    assign n1311 = write[0] ? n287 : \regs[26] [5];   // regs.v(45)
    assign n1312 = write[0] ? n288 : \regs[26] [4];   // regs.v(45)
    assign n1313 = write[0] ? n289 : \regs[26] [3];   // regs.v(45)
    assign n1314 = write[0] ? n290 : \regs[26] [2];   // regs.v(45)
    assign n1315 = write[0] ? n291 : \regs[26] [1];   // regs.v(45)
    assign n1316 = write[0] ? n292 : \regs[26] [0];   // regs.v(45)
    assign n1317 = write[0] ? n293 : \regs[25] [31];   // regs.v(45)
    assign n1318 = write[0] ? n294 : \regs[25] [30];   // regs.v(45)
    assign n1319 = write[0] ? n295 : \regs[25] [29];   // regs.v(45)
    assign n1320 = write[0] ? n296 : \regs[25] [28];   // regs.v(45)
    assign n1321 = write[0] ? n297 : \regs[25] [27];   // regs.v(45)
    assign n1322 = write[0] ? n298 : \regs[25] [26];   // regs.v(45)
    assign n1323 = write[0] ? n299 : \regs[25] [25];   // regs.v(45)
    assign n1324 = write[0] ? n300 : \regs[25] [24];   // regs.v(45)
    assign n1325 = write[0] ? n301 : \regs[25] [23];   // regs.v(45)
    assign n1326 = write[0] ? n302 : \regs[25] [22];   // regs.v(45)
    assign n1327 = write[0] ? n303 : \regs[25] [21];   // regs.v(45)
    assign n1328 = write[0] ? n304 : \regs[25] [20];   // regs.v(45)
    assign n1329 = write[0] ? n305 : \regs[25] [19];   // regs.v(45)
    assign n1330 = write[0] ? n306 : \regs[25] [18];   // regs.v(45)
    assign n1331 = write[0] ? n307 : \regs[25] [17];   // regs.v(45)
    assign n1332 = write[0] ? n308 : \regs[25] [16];   // regs.v(45)
    assign n1333 = write[0] ? n309 : \regs[25] [15];   // regs.v(45)
    assign n1334 = write[0] ? n310 : \regs[25] [14];   // regs.v(45)
    assign n1335 = write[0] ? n311 : \regs[25] [13];   // regs.v(45)
    assign n1336 = write[0] ? n312 : \regs[25] [12];   // regs.v(45)
    assign n1337 = write[0] ? n313 : \regs[25] [11];   // regs.v(45)
    assign n1338 = write[0] ? n314 : \regs[25] [10];   // regs.v(45)
    assign n1339 = write[0] ? n315 : \regs[25] [9];   // regs.v(45)
    assign n1340 = write[0] ? n316 : \regs[25] [8];   // regs.v(45)
    assign n1341 = write[0] ? n317 : \regs[25] [7];   // regs.v(45)
    assign n1342 = write[0] ? n318 : \regs[25] [6];   // regs.v(45)
    assign n1343 = write[0] ? n319 : \regs[25] [5];   // regs.v(45)
    assign n1344 = write[0] ? n320 : \regs[25] [4];   // regs.v(45)
    assign n1345 = write[0] ? n321 : \regs[25] [3];   // regs.v(45)
    assign n1346 = write[0] ? n322 : \regs[25] [2];   // regs.v(45)
    assign n1347 = write[0] ? n323 : \regs[25] [1];   // regs.v(45)
    assign n1348 = write[0] ? n324 : \regs[25] [0];   // regs.v(45)
    assign n1349 = write[0] ? n325 : \regs[24] [31];   // regs.v(45)
    assign n1350 = write[0] ? n326 : \regs[24] [30];   // regs.v(45)
    assign n1351 = write[0] ? n327 : \regs[24] [29];   // regs.v(45)
    assign n1352 = write[0] ? n328 : \regs[24] [28];   // regs.v(45)
    assign n1353 = write[0] ? n329 : \regs[24] [27];   // regs.v(45)
    assign n1354 = write[0] ? n330 : \regs[24] [26];   // regs.v(45)
    assign n1355 = write[0] ? n331 : \regs[24] [25];   // regs.v(45)
    assign n1356 = write[0] ? n332 : \regs[24] [24];   // regs.v(45)
    assign n1357 = write[0] ? n333 : \regs[24] [23];   // regs.v(45)
    assign n1358 = write[0] ? n334 : \regs[24] [22];   // regs.v(45)
    assign n1359 = write[0] ? n335 : \regs[24] [21];   // regs.v(45)
    assign n1360 = write[0] ? n336 : \regs[24] [20];   // regs.v(45)
    assign n1361 = write[0] ? n337 : \regs[24] [19];   // regs.v(45)
    assign n1362 = write[0] ? n338 : \regs[24] [18];   // regs.v(45)
    assign n1363 = write[0] ? n339 : \regs[24] [17];   // regs.v(45)
    assign n1364 = write[0] ? n340 : \regs[24] [16];   // regs.v(45)
    assign n1365 = write[0] ? n341 : \regs[24] [15];   // regs.v(45)
    assign n1366 = write[0] ? n342 : \regs[24] [14];   // regs.v(45)
    assign n1367 = write[0] ? n343 : \regs[24] [13];   // regs.v(45)
    assign n1368 = write[0] ? n344 : \regs[24] [12];   // regs.v(45)
    assign n1369 = write[0] ? n345 : \regs[24] [11];   // regs.v(45)
    assign n1370 = write[0] ? n346 : \regs[24] [10];   // regs.v(45)
    assign n1371 = write[0] ? n347 : \regs[24] [9];   // regs.v(45)
    assign n1372 = write[0] ? n348 : \regs[24] [8];   // regs.v(45)
    assign n1373 = write[0] ? n349 : \regs[24] [7];   // regs.v(45)
    assign n1374 = write[0] ? n350 : \regs[24] [6];   // regs.v(45)
    assign n1375 = write[0] ? n351 : \regs[24] [5];   // regs.v(45)
    assign n1376 = write[0] ? n352 : \regs[24] [4];   // regs.v(45)
    assign n1377 = write[0] ? n353 : \regs[24] [3];   // regs.v(45)
    assign n1378 = write[0] ? n354 : \regs[24] [2];   // regs.v(45)
    assign n1379 = write[0] ? n355 : \regs[24] [1];   // regs.v(45)
    assign n1380 = write[0] ? n356 : \regs[24] [0];   // regs.v(45)
    assign n1381 = write[0] ? n357 : \regs[23] [31];   // regs.v(45)
    assign n1382 = write[0] ? n358 : \regs[23] [30];   // regs.v(45)
    assign n1383 = write[0] ? n359 : \regs[23] [29];   // regs.v(45)
    assign n1384 = write[0] ? n360 : \regs[23] [28];   // regs.v(45)
    assign n1385 = write[0] ? n361 : \regs[23] [27];   // regs.v(45)
    assign n1386 = write[0] ? n362 : \regs[23] [26];   // regs.v(45)
    assign n1387 = write[0] ? n363 : \regs[23] [25];   // regs.v(45)
    assign n1388 = write[0] ? n364 : \regs[23] [24];   // regs.v(45)
    assign n1389 = write[0] ? n365 : \regs[23] [23];   // regs.v(45)
    assign n1390 = write[0] ? n366 : \regs[23] [22];   // regs.v(45)
    assign n1391 = write[0] ? n367 : \regs[23] [21];   // regs.v(45)
    assign n1392 = write[0] ? n368 : \regs[23] [20];   // regs.v(45)
    assign n1393 = write[0] ? n369 : \regs[23] [19];   // regs.v(45)
    assign n1394 = write[0] ? n370 : \regs[23] [18];   // regs.v(45)
    assign n1395 = write[0] ? n371 : \regs[23] [17];   // regs.v(45)
    assign n1396 = write[0] ? n372 : \regs[23] [16];   // regs.v(45)
    assign n1397 = write[0] ? n373 : \regs[23] [15];   // regs.v(45)
    assign n1398 = write[0] ? n374 : \regs[23] [14];   // regs.v(45)
    assign n1399 = write[0] ? n375 : \regs[23] [13];   // regs.v(45)
    assign n1400 = write[0] ? n376 : \regs[23] [12];   // regs.v(45)
    assign n1401 = write[0] ? n377 : \regs[23] [11];   // regs.v(45)
    assign n1402 = write[0] ? n378 : \regs[23] [10];   // regs.v(45)
    assign n1403 = write[0] ? n379 : \regs[23] [9];   // regs.v(45)
    assign n1404 = write[0] ? n380 : \regs[23] [8];   // regs.v(45)
    assign n1405 = write[0] ? n381 : \regs[23] [7];   // regs.v(45)
    assign n1406 = write[0] ? n382 : \regs[23] [6];   // regs.v(45)
    assign n1407 = write[0] ? n383 : \regs[23] [5];   // regs.v(45)
    assign n1408 = write[0] ? n384 : \regs[23] [4];   // regs.v(45)
    assign n1409 = write[0] ? n385 : \regs[23] [3];   // regs.v(45)
    assign n1410 = write[0] ? n386 : \regs[23] [2];   // regs.v(45)
    assign n1411 = write[0] ? n387 : \regs[23] [1];   // regs.v(45)
    assign n1412 = write[0] ? n388 : \regs[23] [0];   // regs.v(45)
    assign n1413 = write[0] ? n389 : \regs[22] [31];   // regs.v(45)
    assign n1414 = write[0] ? n390 : \regs[22] [30];   // regs.v(45)
    assign n1415 = write[0] ? n391 : \regs[22] [29];   // regs.v(45)
    assign n1416 = write[0] ? n392 : \regs[22] [28];   // regs.v(45)
    assign n1417 = write[0] ? n393 : \regs[22] [27];   // regs.v(45)
    assign n1418 = write[0] ? n394 : \regs[22] [26];   // regs.v(45)
    assign n1419 = write[0] ? n395 : \regs[22] [25];   // regs.v(45)
    assign n1420 = write[0] ? n396 : \regs[22] [24];   // regs.v(45)
    assign n1421 = write[0] ? n397 : \regs[22] [23];   // regs.v(45)
    assign n1422 = write[0] ? n398 : \regs[22] [22];   // regs.v(45)
    assign n1423 = write[0] ? n399 : \regs[22] [21];   // regs.v(45)
    assign n1424 = write[0] ? n400 : \regs[22] [20];   // regs.v(45)
    assign n1425 = write[0] ? n401 : \regs[22] [19];   // regs.v(45)
    assign n1426 = write[0] ? n402 : \regs[22] [18];   // regs.v(45)
    assign n1427 = write[0] ? n403 : \regs[22] [17];   // regs.v(45)
    assign n1428 = write[0] ? n404 : \regs[22] [16];   // regs.v(45)
    assign n1429 = write[0] ? n405 : \regs[22] [15];   // regs.v(45)
    assign n1430 = write[0] ? n406 : \regs[22] [14];   // regs.v(45)
    assign n1431 = write[0] ? n407 : \regs[22] [13];   // regs.v(45)
    assign n1432 = write[0] ? n408 : \regs[22] [12];   // regs.v(45)
    assign n1433 = write[0] ? n409 : \regs[22] [11];   // regs.v(45)
    assign n1434 = write[0] ? n410 : \regs[22] [10];   // regs.v(45)
    assign n1435 = write[0] ? n411 : \regs[22] [9];   // regs.v(45)
    assign n1436 = write[0] ? n412 : \regs[22] [8];   // regs.v(45)
    assign n1437 = write[0] ? n413 : \regs[22] [7];   // regs.v(45)
    assign n1438 = write[0] ? n414 : \regs[22] [6];   // regs.v(45)
    assign n1439 = write[0] ? n415 : \regs[22] [5];   // regs.v(45)
    assign n1440 = write[0] ? n416 : \regs[22] [4];   // regs.v(45)
    assign n1441 = write[0] ? n417 : \regs[22] [3];   // regs.v(45)
    assign n1442 = write[0] ? n418 : \regs[22] [2];   // regs.v(45)
    assign n1443 = write[0] ? n419 : \regs[22] [1];   // regs.v(45)
    assign n1444 = write[0] ? n420 : \regs[22] [0];   // regs.v(45)
    assign n1445 = write[0] ? n421 : \regs[21] [31];   // regs.v(45)
    assign n1446 = write[0] ? n422 : \regs[21] [30];   // regs.v(45)
    assign n1447 = write[0] ? n423 : \regs[21] [29];   // regs.v(45)
    assign n1448 = write[0] ? n424 : \regs[21] [28];   // regs.v(45)
    assign n1449 = write[0] ? n425 : \regs[21] [27];   // regs.v(45)
    assign n1450 = write[0] ? n426 : \regs[21] [26];   // regs.v(45)
    assign n1451 = write[0] ? n427 : \regs[21] [25];   // regs.v(45)
    assign n1452 = write[0] ? n428 : \regs[21] [24];   // regs.v(45)
    assign n1453 = write[0] ? n429 : \regs[21] [23];   // regs.v(45)
    assign n1454 = write[0] ? n430 : \regs[21] [22];   // regs.v(45)
    assign n1455 = write[0] ? n431 : \regs[21] [21];   // regs.v(45)
    assign n1456 = write[0] ? n432 : \regs[21] [20];   // regs.v(45)
    assign n1457 = write[0] ? n433 : \regs[21] [19];   // regs.v(45)
    assign n1458 = write[0] ? n434 : \regs[21] [18];   // regs.v(45)
    assign n1459 = write[0] ? n435 : \regs[21] [17];   // regs.v(45)
    assign n1460 = write[0] ? n436 : \regs[21] [16];   // regs.v(45)
    assign n1461 = write[0] ? n437 : \regs[21] [15];   // regs.v(45)
    assign n1462 = write[0] ? n438 : \regs[21] [14];   // regs.v(45)
    assign n1463 = write[0] ? n439 : \regs[21] [13];   // regs.v(45)
    assign n1464 = write[0] ? n440 : \regs[21] [12];   // regs.v(45)
    assign n1465 = write[0] ? n441 : \regs[21] [11];   // regs.v(45)
    assign n1466 = write[0] ? n442 : \regs[21] [10];   // regs.v(45)
    assign n1467 = write[0] ? n443 : \regs[21] [9];   // regs.v(45)
    assign n1468 = write[0] ? n444 : \regs[21] [8];   // regs.v(45)
    assign n1469 = write[0] ? n445 : \regs[21] [7];   // regs.v(45)
    assign n1470 = write[0] ? n446 : \regs[21] [6];   // regs.v(45)
    assign n1471 = write[0] ? n447 : \regs[21] [5];   // regs.v(45)
    assign n1472 = write[0] ? n448 : \regs[21] [4];   // regs.v(45)
    assign n1473 = write[0] ? n449 : \regs[21] [3];   // regs.v(45)
    assign n1474 = write[0] ? n450 : \regs[21] [2];   // regs.v(45)
    assign n1475 = write[0] ? n451 : \regs[21] [1];   // regs.v(45)
    assign n1476 = write[0] ? n452 : \regs[21] [0];   // regs.v(45)
    assign n1477 = write[0] ? n453 : \regs[20] [31];   // regs.v(45)
    assign n1478 = write[0] ? n454 : \regs[20] [30];   // regs.v(45)
    assign n1479 = write[0] ? n455 : \regs[20] [29];   // regs.v(45)
    assign n1480 = write[0] ? n456 : \regs[20] [28];   // regs.v(45)
    assign n1481 = write[0] ? n457 : \regs[20] [27];   // regs.v(45)
    assign n1482 = write[0] ? n458 : \regs[20] [26];   // regs.v(45)
    assign n1483 = write[0] ? n459 : \regs[20] [25];   // regs.v(45)
    assign n1484 = write[0] ? n460 : \regs[20] [24];   // regs.v(45)
    assign n1485 = write[0] ? n461 : \regs[20] [23];   // regs.v(45)
    assign n1486 = write[0] ? n462 : \regs[20] [22];   // regs.v(45)
    assign n1487 = write[0] ? n463 : \regs[20] [21];   // regs.v(45)
    assign n1488 = write[0] ? n464 : \regs[20] [20];   // regs.v(45)
    assign n1489 = write[0] ? n465 : \regs[20] [19];   // regs.v(45)
    assign n1490 = write[0] ? n466 : \regs[20] [18];   // regs.v(45)
    assign n1491 = write[0] ? n467 : \regs[20] [17];   // regs.v(45)
    assign n1492 = write[0] ? n468 : \regs[20] [16];   // regs.v(45)
    assign n1493 = write[0] ? n469 : \regs[20] [15];   // regs.v(45)
    assign n1494 = write[0] ? n470 : \regs[20] [14];   // regs.v(45)
    assign n1495 = write[0] ? n471 : \regs[20] [13];   // regs.v(45)
    assign n1496 = write[0] ? n472 : \regs[20] [12];   // regs.v(45)
    assign n1497 = write[0] ? n473 : \regs[20] [11];   // regs.v(45)
    assign n1498 = write[0] ? n474 : \regs[20] [10];   // regs.v(45)
    assign n1499 = write[0] ? n475 : \regs[20] [9];   // regs.v(45)
    assign n1500 = write[0] ? n476 : \regs[20] [8];   // regs.v(45)
    assign n1501 = write[0] ? n477 : \regs[20] [7];   // regs.v(45)
    assign n1502 = write[0] ? n478 : \regs[20] [6];   // regs.v(45)
    assign n1503 = write[0] ? n479 : \regs[20] [5];   // regs.v(45)
    assign n1504 = write[0] ? n480 : \regs[20] [4];   // regs.v(45)
    assign n1505 = write[0] ? n481 : \regs[20] [3];   // regs.v(45)
    assign n1506 = write[0] ? n482 : \regs[20] [2];   // regs.v(45)
    assign n1507 = write[0] ? n483 : \regs[20] [1];   // regs.v(45)
    assign n1508 = write[0] ? n484 : \regs[20] [0];   // regs.v(45)
    assign n1509 = write[0] ? n485 : \regs[19] [31];   // regs.v(45)
    assign n1510 = write[0] ? n486 : \regs[19] [30];   // regs.v(45)
    assign n1511 = write[0] ? n487 : \regs[19] [29];   // regs.v(45)
    assign n1512 = write[0] ? n488 : \regs[19] [28];   // regs.v(45)
    assign n1513 = write[0] ? n489 : \regs[19] [27];   // regs.v(45)
    assign n1514 = write[0] ? n490 : \regs[19] [26];   // regs.v(45)
    assign n1515 = write[0] ? n491 : \regs[19] [25];   // regs.v(45)
    assign n1516 = write[0] ? n492 : \regs[19] [24];   // regs.v(45)
    assign n1517 = write[0] ? n493 : \regs[19] [23];   // regs.v(45)
    assign n1518 = write[0] ? n494 : \regs[19] [22];   // regs.v(45)
    assign n1519 = write[0] ? n495 : \regs[19] [21];   // regs.v(45)
    assign n1520 = write[0] ? n496 : \regs[19] [20];   // regs.v(45)
    assign n1521 = write[0] ? n497 : \regs[19] [19];   // regs.v(45)
    assign n1522 = write[0] ? n498 : \regs[19] [18];   // regs.v(45)
    assign n1523 = write[0] ? n499 : \regs[19] [17];   // regs.v(45)
    assign n1524 = write[0] ? n500 : \regs[19] [16];   // regs.v(45)
    assign n1525 = write[0] ? n501 : \regs[19] [15];   // regs.v(45)
    assign n1526 = write[0] ? n502 : \regs[19] [14];   // regs.v(45)
    assign n1527 = write[0] ? n503 : \regs[19] [13];   // regs.v(45)
    assign n1528 = write[0] ? n504 : \regs[19] [12];   // regs.v(45)
    assign n1529 = write[0] ? n505 : \regs[19] [11];   // regs.v(45)
    assign n1530 = write[0] ? n506 : \regs[19] [10];   // regs.v(45)
    assign n1531 = write[0] ? n507 : \regs[19] [9];   // regs.v(45)
    assign n1532 = write[0] ? n508 : \regs[19] [8];   // regs.v(45)
    assign n1533 = write[0] ? n509 : \regs[19] [7];   // regs.v(45)
    assign n1534 = write[0] ? n510 : \regs[19] [6];   // regs.v(45)
    assign n1535 = write[0] ? n511 : \regs[19] [5];   // regs.v(45)
    assign n1536 = write[0] ? n512 : \regs[19] [4];   // regs.v(45)
    assign n1537 = write[0] ? n513 : \regs[19] [3];   // regs.v(45)
    assign n1538 = write[0] ? n514 : \regs[19] [2];   // regs.v(45)
    assign n1539 = write[0] ? n515 : \regs[19] [1];   // regs.v(45)
    assign n1540 = write[0] ? n516 : \regs[19] [0];   // regs.v(45)
    assign n1541 = write[0] ? n517 : \regs[18] [31];   // regs.v(45)
    assign n1542 = write[0] ? n518 : \regs[18] [30];   // regs.v(45)
    assign n1543 = write[0] ? n519 : \regs[18] [29];   // regs.v(45)
    assign n1544 = write[0] ? n520 : \regs[18] [28];   // regs.v(45)
    assign n1545 = write[0] ? n521 : \regs[18] [27];   // regs.v(45)
    assign n1546 = write[0] ? n522 : \regs[18] [26];   // regs.v(45)
    assign n1547 = write[0] ? n523 : \regs[18] [25];   // regs.v(45)
    assign n1548 = write[0] ? n524 : \regs[18] [24];   // regs.v(45)
    assign n1549 = write[0] ? n525 : \regs[18] [23];   // regs.v(45)
    assign n1550 = write[0] ? n526 : \regs[18] [22];   // regs.v(45)
    assign n1551 = write[0] ? n527 : \regs[18] [21];   // regs.v(45)
    assign n1552 = write[0] ? n528 : \regs[18] [20];   // regs.v(45)
    assign n1553 = write[0] ? n529 : \regs[18] [19];   // regs.v(45)
    assign n1554 = write[0] ? n530 : \regs[18] [18];   // regs.v(45)
    assign n1555 = write[0] ? n531 : \regs[18] [17];   // regs.v(45)
    assign n1556 = write[0] ? n532 : \regs[18] [16];   // regs.v(45)
    assign n1557 = write[0] ? n533 : \regs[18] [15];   // regs.v(45)
    assign n1558 = write[0] ? n534 : \regs[18] [14];   // regs.v(45)
    assign n1559 = write[0] ? n535 : \regs[18] [13];   // regs.v(45)
    assign n1560 = write[0] ? n536 : \regs[18] [12];   // regs.v(45)
    assign n1561 = write[0] ? n537 : \regs[18] [11];   // regs.v(45)
    assign n1562 = write[0] ? n538 : \regs[18] [10];   // regs.v(45)
    assign n1563 = write[0] ? n539 : \regs[18] [9];   // regs.v(45)
    assign n1564 = write[0] ? n540 : \regs[18] [8];   // regs.v(45)
    assign n1565 = write[0] ? n541 : \regs[18] [7];   // regs.v(45)
    assign n1566 = write[0] ? n542 : \regs[18] [6];   // regs.v(45)
    assign n1567 = write[0] ? n543 : \regs[18] [5];   // regs.v(45)
    assign n1568 = write[0] ? n544 : \regs[18] [4];   // regs.v(45)
    assign n1569 = write[0] ? n545 : \regs[18] [3];   // regs.v(45)
    assign n1570 = write[0] ? n546 : \regs[18] [2];   // regs.v(45)
    assign n1571 = write[0] ? n547 : \regs[18] [1];   // regs.v(45)
    assign n1572 = write[0] ? n548 : \regs[18] [0];   // regs.v(45)
    assign n1573 = write[0] ? n549 : \regs[17] [31];   // regs.v(45)
    assign n1574 = write[0] ? n550 : \regs[17] [30];   // regs.v(45)
    assign n1575 = write[0] ? n551 : \regs[17] [29];   // regs.v(45)
    assign n1576 = write[0] ? n552 : \regs[17] [28];   // regs.v(45)
    assign n1577 = write[0] ? n553 : \regs[17] [27];   // regs.v(45)
    assign n1578 = write[0] ? n554 : \regs[17] [26];   // regs.v(45)
    assign n1579 = write[0] ? n555 : \regs[17] [25];   // regs.v(45)
    assign n1580 = write[0] ? n556 : \regs[17] [24];   // regs.v(45)
    assign n1581 = write[0] ? n557 : \regs[17] [23];   // regs.v(45)
    assign n1582 = write[0] ? n558 : \regs[17] [22];   // regs.v(45)
    assign n1583 = write[0] ? n559 : \regs[17] [21];   // regs.v(45)
    assign n1584 = write[0] ? n560 : \regs[17] [20];   // regs.v(45)
    assign n1585 = write[0] ? n561 : \regs[17] [19];   // regs.v(45)
    assign n1586 = write[0] ? n562 : \regs[17] [18];   // regs.v(45)
    assign n1587 = write[0] ? n563 : \regs[17] [17];   // regs.v(45)
    assign n1588 = write[0] ? n564 : \regs[17] [16];   // regs.v(45)
    assign n1589 = write[0] ? n565 : \regs[17] [15];   // regs.v(45)
    assign n1590 = write[0] ? n566 : \regs[17] [14];   // regs.v(45)
    assign n1591 = write[0] ? n567 : \regs[17] [13];   // regs.v(45)
    assign n1592 = write[0] ? n568 : \regs[17] [12];   // regs.v(45)
    assign n1593 = write[0] ? n569 : \regs[17] [11];   // regs.v(45)
    assign n1594 = write[0] ? n570 : \regs[17] [10];   // regs.v(45)
    assign n1595 = write[0] ? n571 : \regs[17] [9];   // regs.v(45)
    assign n1596 = write[0] ? n572 : \regs[17] [8];   // regs.v(45)
    assign n1597 = write[0] ? n573 : \regs[17] [7];   // regs.v(45)
    assign n1598 = write[0] ? n574 : \regs[17] [6];   // regs.v(45)
    assign n1599 = write[0] ? n575 : \regs[17] [5];   // regs.v(45)
    assign n1600 = write[0] ? n576 : \regs[17] [4];   // regs.v(45)
    assign n1601 = write[0] ? n577 : \regs[17] [3];   // regs.v(45)
    assign n1602 = write[0] ? n578 : \regs[17] [2];   // regs.v(45)
    assign n1603 = write[0] ? n579 : \regs[17] [1];   // regs.v(45)
    assign n1604 = write[0] ? n580 : \regs[17] [0];   // regs.v(45)
    assign n1605 = write[0] ? n581 : \regs[16] [31];   // regs.v(45)
    assign n1606 = write[0] ? n582 : \regs[16] [30];   // regs.v(45)
    assign n1607 = write[0] ? n583 : \regs[16] [29];   // regs.v(45)
    assign n1608 = write[0] ? n584 : \regs[16] [28];   // regs.v(45)
    assign n1609 = write[0] ? n585 : \regs[16] [27];   // regs.v(45)
    assign n1610 = write[0] ? n586 : \regs[16] [26];   // regs.v(45)
    assign n1611 = write[0] ? n587 : \regs[16] [25];   // regs.v(45)
    assign n1612 = write[0] ? n588 : \regs[16] [24];   // regs.v(45)
    assign n1613 = write[0] ? n589 : \regs[16] [23];   // regs.v(45)
    assign n1614 = write[0] ? n590 : \regs[16] [22];   // regs.v(45)
    assign n1615 = write[0] ? n591 : \regs[16] [21];   // regs.v(45)
    assign n1616 = write[0] ? n592 : \regs[16] [20];   // regs.v(45)
    assign n1617 = write[0] ? n593 : \regs[16] [19];   // regs.v(45)
    assign n1618 = write[0] ? n594 : \regs[16] [18];   // regs.v(45)
    assign n1619 = write[0] ? n595 : \regs[16] [17];   // regs.v(45)
    assign n1620 = write[0] ? n596 : \regs[16] [16];   // regs.v(45)
    assign n1621 = write[0] ? n597 : \regs[16] [15];   // regs.v(45)
    assign n1622 = write[0] ? n598 : \regs[16] [14];   // regs.v(45)
    assign n1623 = write[0] ? n599 : \regs[16] [13];   // regs.v(45)
    assign n1624 = write[0] ? n600 : \regs[16] [12];   // regs.v(45)
    assign n1625 = write[0] ? n601 : \regs[16] [11];   // regs.v(45)
    assign n1626 = write[0] ? n602 : \regs[16] [10];   // regs.v(45)
    assign n1627 = write[0] ? n603 : \regs[16] [9];   // regs.v(45)
    assign n1628 = write[0] ? n604 : \regs[16] [8];   // regs.v(45)
    assign n1629 = write[0] ? n605 : \regs[16] [7];   // regs.v(45)
    assign n1630 = write[0] ? n606 : \regs[16] [6];   // regs.v(45)
    assign n1631 = write[0] ? n607 : \regs[16] [5];   // regs.v(45)
    assign n1632 = write[0] ? n608 : \regs[16] [4];   // regs.v(45)
    assign n1633 = write[0] ? n609 : \regs[16] [3];   // regs.v(45)
    assign n1634 = write[0] ? n610 : \regs[16] [2];   // regs.v(45)
    assign n1635 = write[0] ? n611 : \regs[16] [1];   // regs.v(45)
    assign n1636 = write[0] ? n612 : \regs[16] [0];   // regs.v(45)
    assign n1637 = write[0] ? n613 : \regs[15] [31];   // regs.v(45)
    assign n1638 = write[0] ? n614 : \regs[15] [30];   // regs.v(45)
    assign n1639 = write[0] ? n615 : \regs[15] [29];   // regs.v(45)
    assign n1640 = write[0] ? n616 : \regs[15] [28];   // regs.v(45)
    assign n1641 = write[0] ? n617 : \regs[15] [27];   // regs.v(45)
    assign n1642 = write[0] ? n618 : \regs[15] [26];   // regs.v(45)
    assign n1643 = write[0] ? n619 : \regs[15] [25];   // regs.v(45)
    assign n1644 = write[0] ? n620 : \regs[15] [24];   // regs.v(45)
    assign n1645 = write[0] ? n621 : \regs[15] [23];   // regs.v(45)
    assign n1646 = write[0] ? n622 : \regs[15] [22];   // regs.v(45)
    assign n1647 = write[0] ? n623 : \regs[15] [21];   // regs.v(45)
    assign n1648 = write[0] ? n624 : \regs[15] [20];   // regs.v(45)
    assign n1649 = write[0] ? n625 : \regs[15] [19];   // regs.v(45)
    assign n1650 = write[0] ? n626 : \regs[15] [18];   // regs.v(45)
    assign n1651 = write[0] ? n627 : \regs[15] [17];   // regs.v(45)
    assign n1652 = write[0] ? n628 : \regs[15] [16];   // regs.v(45)
    assign n1653 = write[0] ? n629 : \regs[15] [15];   // regs.v(45)
    assign n1654 = write[0] ? n630 : \regs[15] [14];   // regs.v(45)
    assign n1655 = write[0] ? n631 : \regs[15] [13];   // regs.v(45)
    assign n1656 = write[0] ? n632 : \regs[15] [12];   // regs.v(45)
    assign n1657 = write[0] ? n633 : \regs[15] [11];   // regs.v(45)
    assign n1658 = write[0] ? n634 : \regs[15] [10];   // regs.v(45)
    assign n1659 = write[0] ? n635 : \regs[15] [9];   // regs.v(45)
    assign n1660 = write[0] ? n636 : \regs[15] [8];   // regs.v(45)
    assign n1661 = write[0] ? n637 : \regs[15] [7];   // regs.v(45)
    assign n1662 = write[0] ? n638 : \regs[15] [6];   // regs.v(45)
    assign n1663 = write[0] ? n639 : \regs[15] [5];   // regs.v(45)
    assign n1664 = write[0] ? n640 : \regs[15] [4];   // regs.v(45)
    assign n1665 = write[0] ? n641 : \regs[15] [3];   // regs.v(45)
    assign n1666 = write[0] ? n642 : \regs[15] [2];   // regs.v(45)
    assign n1667 = write[0] ? n643 : \regs[15] [1];   // regs.v(45)
    assign n1668 = write[0] ? n644 : \regs[15] [0];   // regs.v(45)
    assign n1669 = write[0] ? n645 : \regs[14] [31];   // regs.v(45)
    assign n1670 = write[0] ? n646 : \regs[14] [30];   // regs.v(45)
    assign n1671 = write[0] ? n647 : \regs[14] [29];   // regs.v(45)
    assign n1672 = write[0] ? n648 : \regs[14] [28];   // regs.v(45)
    assign n1673 = write[0] ? n649 : \regs[14] [27];   // regs.v(45)
    assign n1674 = write[0] ? n650 : \regs[14] [26];   // regs.v(45)
    assign n1675 = write[0] ? n651 : \regs[14] [25];   // regs.v(45)
    assign n1676 = write[0] ? n652 : \regs[14] [24];   // regs.v(45)
    assign n1677 = write[0] ? n653 : \regs[14] [23];   // regs.v(45)
    assign n1678 = write[0] ? n654 : \regs[14] [22];   // regs.v(45)
    assign n1679 = write[0] ? n655 : \regs[14] [21];   // regs.v(45)
    assign n1680 = write[0] ? n656 : \regs[14] [20];   // regs.v(45)
    assign n1681 = write[0] ? n657 : \regs[14] [19];   // regs.v(45)
    assign n1682 = write[0] ? n658 : \regs[14] [18];   // regs.v(45)
    assign n1683 = write[0] ? n659 : \regs[14] [17];   // regs.v(45)
    assign n1684 = write[0] ? n660 : \regs[14] [16];   // regs.v(45)
    assign n1685 = write[0] ? n661 : \regs[14] [15];   // regs.v(45)
    assign n1686 = write[0] ? n662 : \regs[14] [14];   // regs.v(45)
    assign n1687 = write[0] ? n663 : \regs[14] [13];   // regs.v(45)
    assign n1688 = write[0] ? n664 : \regs[14] [12];   // regs.v(45)
    assign n1689 = write[0] ? n665 : \regs[14] [11];   // regs.v(45)
    assign n1690 = write[0] ? n666 : \regs[14] [10];   // regs.v(45)
    assign n1691 = write[0] ? n667 : \regs[14] [9];   // regs.v(45)
    assign n1692 = write[0] ? n668 : \regs[14] [8];   // regs.v(45)
    assign n1693 = write[0] ? n669 : \regs[14] [7];   // regs.v(45)
    assign n1694 = write[0] ? n670 : \regs[14] [6];   // regs.v(45)
    assign n1695 = write[0] ? n671 : \regs[14] [5];   // regs.v(45)
    assign n1696 = write[0] ? n672 : \regs[14] [4];   // regs.v(45)
    assign n1697 = write[0] ? n673 : \regs[14] [3];   // regs.v(45)
    assign n1698 = write[0] ? n674 : \regs[14] [2];   // regs.v(45)
    assign n1699 = write[0] ? n675 : \regs[14] [1];   // regs.v(45)
    assign n1700 = write[0] ? n676 : \regs[14] [0];   // regs.v(45)
    assign n1701 = write[0] ? n677 : \regs[13] [31];   // regs.v(45)
    assign n1702 = write[0] ? n678 : \regs[13] [30];   // regs.v(45)
    assign n1703 = write[0] ? n679 : \regs[13] [29];   // regs.v(45)
    assign n1704 = write[0] ? n680 : \regs[13] [28];   // regs.v(45)
    assign n1705 = write[0] ? n681 : \regs[13] [27];   // regs.v(45)
    assign n1706 = write[0] ? n682 : \regs[13] [26];   // regs.v(45)
    assign n1707 = write[0] ? n683 : \regs[13] [25];   // regs.v(45)
    assign n1708 = write[0] ? n684 : \regs[13] [24];   // regs.v(45)
    assign n1709 = write[0] ? n685 : \regs[13] [23];   // regs.v(45)
    assign n1710 = write[0] ? n686 : \regs[13] [22];   // regs.v(45)
    assign n1711 = write[0] ? n687 : \regs[13] [21];   // regs.v(45)
    assign n1712 = write[0] ? n688 : \regs[13] [20];   // regs.v(45)
    assign n1713 = write[0] ? n689 : \regs[13] [19];   // regs.v(45)
    assign n1714 = write[0] ? n690 : \regs[13] [18];   // regs.v(45)
    assign n1715 = write[0] ? n691 : \regs[13] [17];   // regs.v(45)
    assign n1716 = write[0] ? n692 : \regs[13] [16];   // regs.v(45)
    assign n1717 = write[0] ? n693 : \regs[13] [15];   // regs.v(45)
    assign n1718 = write[0] ? n694 : \regs[13] [14];   // regs.v(45)
    assign n1719 = write[0] ? n695 : \regs[13] [13];   // regs.v(45)
    assign n1720 = write[0] ? n696 : \regs[13] [12];   // regs.v(45)
    assign n1721 = write[0] ? n697 : \regs[13] [11];   // regs.v(45)
    assign n1722 = write[0] ? n698 : \regs[13] [10];   // regs.v(45)
    assign n1723 = write[0] ? n699 : \regs[13] [9];   // regs.v(45)
    assign n1724 = write[0] ? n700 : \regs[13] [8];   // regs.v(45)
    assign n1725 = write[0] ? n701 : \regs[13] [7];   // regs.v(45)
    assign n1726 = write[0] ? n702 : \regs[13] [6];   // regs.v(45)
    assign n1727 = write[0] ? n703 : \regs[13] [5];   // regs.v(45)
    assign n1728 = write[0] ? n704 : \regs[13] [4];   // regs.v(45)
    assign n1729 = write[0] ? n705 : \regs[13] [3];   // regs.v(45)
    assign n1730 = write[0] ? n706 : \regs[13] [2];   // regs.v(45)
    assign n1731 = write[0] ? n707 : \regs[13] [1];   // regs.v(45)
    assign n1732 = write[0] ? n708 : \regs[13] [0];   // regs.v(45)
    assign n1733 = write[0] ? n709 : \regs[12] [31];   // regs.v(45)
    assign n1734 = write[0] ? n710 : \regs[12] [30];   // regs.v(45)
    assign n1735 = write[0] ? n711 : \regs[12] [29];   // regs.v(45)
    assign n1736 = write[0] ? n712 : \regs[12] [28];   // regs.v(45)
    assign n1737 = write[0] ? n713 : \regs[12] [27];   // regs.v(45)
    assign n1738 = write[0] ? n714 : \regs[12] [26];   // regs.v(45)
    assign n1739 = write[0] ? n715 : \regs[12] [25];   // regs.v(45)
    assign n1740 = write[0] ? n716 : \regs[12] [24];   // regs.v(45)
    assign n1741 = write[0] ? n717 : \regs[12] [23];   // regs.v(45)
    assign n1742 = write[0] ? n718 : \regs[12] [22];   // regs.v(45)
    assign n1743 = write[0] ? n719 : \regs[12] [21];   // regs.v(45)
    assign n1744 = write[0] ? n720 : \regs[12] [20];   // regs.v(45)
    assign n1745 = write[0] ? n721 : \regs[12] [19];   // regs.v(45)
    assign n1746 = write[0] ? n722 : \regs[12] [18];   // regs.v(45)
    assign n1747 = write[0] ? n723 : \regs[12] [17];   // regs.v(45)
    assign n1748 = write[0] ? n724 : \regs[12] [16];   // regs.v(45)
    assign n1749 = write[0] ? n725 : \regs[12] [15];   // regs.v(45)
    assign n1750 = write[0] ? n726 : \regs[12] [14];   // regs.v(45)
    assign n1751 = write[0] ? n727 : \regs[12] [13];   // regs.v(45)
    assign n1752 = write[0] ? n728 : \regs[12] [12];   // regs.v(45)
    assign n1753 = write[0] ? n729 : \regs[12] [11];   // regs.v(45)
    assign n1754 = write[0] ? n730 : \regs[12] [10];   // regs.v(45)
    assign n1755 = write[0] ? n731 : \regs[12] [9];   // regs.v(45)
    assign n1756 = write[0] ? n732 : \regs[12] [8];   // regs.v(45)
    assign n1757 = write[0] ? n733 : \regs[12] [7];   // regs.v(45)
    assign n1758 = write[0] ? n734 : \regs[12] [6];   // regs.v(45)
    assign n1759 = write[0] ? n735 : \regs[12] [5];   // regs.v(45)
    assign n1760 = write[0] ? n736 : \regs[12] [4];   // regs.v(45)
    assign n1761 = write[0] ? n737 : \regs[12] [3];   // regs.v(45)
    assign n1762 = write[0] ? n738 : \regs[12] [2];   // regs.v(45)
    assign n1763 = write[0] ? n739 : \regs[12] [1];   // regs.v(45)
    assign n1764 = write[0] ? n740 : \regs[12] [0];   // regs.v(45)
    assign n1765 = write[0] ? n741 : \regs[11] [31];   // regs.v(45)
    assign n1766 = write[0] ? n742 : \regs[11] [30];   // regs.v(45)
    assign n1767 = write[0] ? n743 : \regs[11] [29];   // regs.v(45)
    assign n1768 = write[0] ? n744 : \regs[11] [28];   // regs.v(45)
    assign n1769 = write[0] ? n745 : \regs[11] [27];   // regs.v(45)
    assign n1770 = write[0] ? n746 : \regs[11] [26];   // regs.v(45)
    assign n1771 = write[0] ? n747 : \regs[11] [25];   // regs.v(45)
    assign n1772 = write[0] ? n748 : \regs[11] [24];   // regs.v(45)
    assign n1773 = write[0] ? n749 : \regs[11] [23];   // regs.v(45)
    assign n1774 = write[0] ? n750 : \regs[11] [22];   // regs.v(45)
    assign n1775 = write[0] ? n751 : \regs[11] [21];   // regs.v(45)
    assign n1776 = write[0] ? n752 : \regs[11] [20];   // regs.v(45)
    assign n1777 = write[0] ? n753 : \regs[11] [19];   // regs.v(45)
    assign n1778 = write[0] ? n754 : \regs[11] [18];   // regs.v(45)
    assign n1779 = write[0] ? n755 : \regs[11] [17];   // regs.v(45)
    assign n1780 = write[0] ? n756 : \regs[11] [16];   // regs.v(45)
    assign n1781 = write[0] ? n757 : \regs[11] [15];   // regs.v(45)
    assign n1782 = write[0] ? n758 : \regs[11] [14];   // regs.v(45)
    assign n1783 = write[0] ? n759 : \regs[11] [13];   // regs.v(45)
    assign n1784 = write[0] ? n760 : \regs[11] [12];   // regs.v(45)
    assign n1785 = write[0] ? n761 : \regs[11] [11];   // regs.v(45)
    assign n1786 = write[0] ? n762 : \regs[11] [10];   // regs.v(45)
    assign n1787 = write[0] ? n763 : \regs[11] [9];   // regs.v(45)
    assign n1788 = write[0] ? n764 : \regs[11] [8];   // regs.v(45)
    assign n1789 = write[0] ? n765 : \regs[11] [7];   // regs.v(45)
    assign n1790 = write[0] ? n766 : \regs[11] [6];   // regs.v(45)
    assign n1791 = write[0] ? n767 : \regs[11] [5];   // regs.v(45)
    assign n1792 = write[0] ? n768 : \regs[11] [4];   // regs.v(45)
    assign n1793 = write[0] ? n769 : \regs[11] [3];   // regs.v(45)
    assign n1794 = write[0] ? n770 : \regs[11] [2];   // regs.v(45)
    assign n1795 = write[0] ? n771 : \regs[11] [1];   // regs.v(45)
    assign n1796 = write[0] ? n772 : \regs[11] [0];   // regs.v(45)
    assign n1797 = write[0] ? n773 : \regs[10] [31];   // regs.v(45)
    assign n1798 = write[0] ? n774 : \regs[10] [30];   // regs.v(45)
    assign n1799 = write[0] ? n775 : \regs[10] [29];   // regs.v(45)
    assign n1800 = write[0] ? n776 : \regs[10] [28];   // regs.v(45)
    assign n1801 = write[0] ? n777 : \regs[10] [27];   // regs.v(45)
    assign n1802 = write[0] ? n778 : \regs[10] [26];   // regs.v(45)
    assign n1803 = write[0] ? n779 : \regs[10] [25];   // regs.v(45)
    assign n1804 = write[0] ? n780 : \regs[10] [24];   // regs.v(45)
    assign n1805 = write[0] ? n781 : \regs[10] [23];   // regs.v(45)
    assign n1806 = write[0] ? n782 : \regs[10] [22];   // regs.v(45)
    assign n1807 = write[0] ? n783 : \regs[10] [21];   // regs.v(45)
    assign n1808 = write[0] ? n784 : \regs[10] [20];   // regs.v(45)
    assign n1809 = write[0] ? n785 : \regs[10] [19];   // regs.v(45)
    assign n1810 = write[0] ? n786 : \regs[10] [18];   // regs.v(45)
    assign n1811 = write[0] ? n787 : \regs[10] [17];   // regs.v(45)
    assign n1812 = write[0] ? n788 : \regs[10] [16];   // regs.v(45)
    assign n1813 = write[0] ? n789 : \regs[10] [15];   // regs.v(45)
    assign n1814 = write[0] ? n790 : \regs[10] [14];   // regs.v(45)
    assign n1815 = write[0] ? n791 : \regs[10] [13];   // regs.v(45)
    assign n1816 = write[0] ? n792 : \regs[10] [12];   // regs.v(45)
    assign n1817 = write[0] ? n793 : \regs[10] [11];   // regs.v(45)
    assign n1818 = write[0] ? n794 : \regs[10] [10];   // regs.v(45)
    assign n1819 = write[0] ? n795 : \regs[10] [9];   // regs.v(45)
    assign n1820 = write[0] ? n796 : \regs[10] [8];   // regs.v(45)
    assign n1821 = write[0] ? n797 : \regs[10] [7];   // regs.v(45)
    assign n1822 = write[0] ? n798 : \regs[10] [6];   // regs.v(45)
    assign n1823 = write[0] ? n799 : \regs[10] [5];   // regs.v(45)
    assign n1824 = write[0] ? n800 : \regs[10] [4];   // regs.v(45)
    assign n1825 = write[0] ? n801 : \regs[10] [3];   // regs.v(45)
    assign n1826 = write[0] ? n802 : \regs[10] [2];   // regs.v(45)
    assign n1827 = write[0] ? n803 : \regs[10] [1];   // regs.v(45)
    assign n1828 = write[0] ? n804 : \regs[10] [0];   // regs.v(45)
    assign n1829 = write[0] ? n805 : \regs[9] [31];   // regs.v(45)
    assign n1830 = write[0] ? n806 : \regs[9] [30];   // regs.v(45)
    assign n1831 = write[0] ? n807 : \regs[9] [29];   // regs.v(45)
    assign n1832 = write[0] ? n808 : \regs[9] [28];   // regs.v(45)
    assign n1833 = write[0] ? n809 : \regs[9] [27];   // regs.v(45)
    assign n1834 = write[0] ? n810 : \regs[9] [26];   // regs.v(45)
    assign n1835 = write[0] ? n811 : \regs[9] [25];   // regs.v(45)
    assign n1836 = write[0] ? n812 : \regs[9] [24];   // regs.v(45)
    assign n1837 = write[0] ? n813 : \regs[9] [23];   // regs.v(45)
    assign n1838 = write[0] ? n814 : \regs[9] [22];   // regs.v(45)
    assign n1839 = write[0] ? n815 : \regs[9] [21];   // regs.v(45)
    assign n1840 = write[0] ? n816 : \regs[9] [20];   // regs.v(45)
    assign n1841 = write[0] ? n817 : \regs[9] [19];   // regs.v(45)
    assign n1842 = write[0] ? n818 : \regs[9] [18];   // regs.v(45)
    assign n1843 = write[0] ? n819 : \regs[9] [17];   // regs.v(45)
    assign n1844 = write[0] ? n820 : \regs[9] [16];   // regs.v(45)
    assign n1845 = write[0] ? n821 : \regs[9] [15];   // regs.v(45)
    assign n1846 = write[0] ? n822 : \regs[9] [14];   // regs.v(45)
    assign n1847 = write[0] ? n823 : \regs[9] [13];   // regs.v(45)
    assign n1848 = write[0] ? n824 : \regs[9] [12];   // regs.v(45)
    assign n1849 = write[0] ? n825 : \regs[9] [11];   // regs.v(45)
    assign n1850 = write[0] ? n826 : \regs[9] [10];   // regs.v(45)
    assign n1851 = write[0] ? n827 : \regs[9] [9];   // regs.v(45)
    assign n1852 = write[0] ? n828 : \regs[9] [8];   // regs.v(45)
    assign n1853 = write[0] ? n829 : \regs[9] [7];   // regs.v(45)
    assign n1854 = write[0] ? n830 : \regs[9] [6];   // regs.v(45)
    assign n1855 = write[0] ? n831 : \regs[9] [5];   // regs.v(45)
    assign n1856 = write[0] ? n832 : \regs[9] [4];   // regs.v(45)
    assign n1857 = write[0] ? n833 : \regs[9] [3];   // regs.v(45)
    assign n1858 = write[0] ? n834 : \regs[9] [2];   // regs.v(45)
    assign n1859 = write[0] ? n835 : \regs[9] [1];   // regs.v(45)
    assign n1860 = write[0] ? n836 : \regs[9] [0];   // regs.v(45)
    assign n1861 = write[0] ? n837 : \regs[8] [31];   // regs.v(45)
    assign n1862 = write[0] ? n838 : \regs[8] [30];   // regs.v(45)
    assign n1863 = write[0] ? n839 : \regs[8] [29];   // regs.v(45)
    assign n1864 = write[0] ? n840 : \regs[8] [28];   // regs.v(45)
    assign n1865 = write[0] ? n841 : \regs[8] [27];   // regs.v(45)
    assign n1866 = write[0] ? n842 : \regs[8] [26];   // regs.v(45)
    assign n1867 = write[0] ? n843 : \regs[8] [25];   // regs.v(45)
    assign n1868 = write[0] ? n844 : \regs[8] [24];   // regs.v(45)
    assign n1869 = write[0] ? n845 : \regs[8] [23];   // regs.v(45)
    assign n1870 = write[0] ? n846 : \regs[8] [22];   // regs.v(45)
    assign n1871 = write[0] ? n847 : \regs[8] [21];   // regs.v(45)
    assign n1872 = write[0] ? n848 : \regs[8] [20];   // regs.v(45)
    assign n1873 = write[0] ? n849 : \regs[8] [19];   // regs.v(45)
    assign n1874 = write[0] ? n850 : \regs[8] [18];   // regs.v(45)
    assign n1875 = write[0] ? n851 : \regs[8] [17];   // regs.v(45)
    assign n1876 = write[0] ? n852 : \regs[8] [16];   // regs.v(45)
    assign n1877 = write[0] ? n853 : \regs[8] [15];   // regs.v(45)
    assign n1878 = write[0] ? n854 : \regs[8] [14];   // regs.v(45)
    assign n1879 = write[0] ? n855 : \regs[8] [13];   // regs.v(45)
    assign n1880 = write[0] ? n856 : \regs[8] [12];   // regs.v(45)
    assign n1881 = write[0] ? n857 : \regs[8] [11];   // regs.v(45)
    assign n1882 = write[0] ? n858 : \regs[8] [10];   // regs.v(45)
    assign n1883 = write[0] ? n859 : \regs[8] [9];   // regs.v(45)
    assign n1884 = write[0] ? n860 : \regs[8] [8];   // regs.v(45)
    assign n1885 = write[0] ? n861 : \regs[8] [7];   // regs.v(45)
    assign n1886 = write[0] ? n862 : \regs[8] [6];   // regs.v(45)
    assign n1887 = write[0] ? n863 : \regs[8] [5];   // regs.v(45)
    assign n1888 = write[0] ? n864 : \regs[8] [4];   // regs.v(45)
    assign n1889 = write[0] ? n865 : \regs[8] [3];   // regs.v(45)
    assign n1890 = write[0] ? n866 : \regs[8] [2];   // regs.v(45)
    assign n1891 = write[0] ? n867 : \regs[8] [1];   // regs.v(45)
    assign n1892 = write[0] ? n868 : \regs[8] [0];   // regs.v(45)
    assign n1893 = write[0] ? n869 : \regs[7] [31];   // regs.v(45)
    assign n1894 = write[0] ? n870 : \regs[7] [30];   // regs.v(45)
    assign n1895 = write[0] ? n871 : \regs[7] [29];   // regs.v(45)
    assign n1896 = write[0] ? n872 : \regs[7] [28];   // regs.v(45)
    assign n1897 = write[0] ? n873 : \regs[7] [27];   // regs.v(45)
    assign n1898 = write[0] ? n874 : \regs[7] [26];   // regs.v(45)
    assign n1899 = write[0] ? n875 : \regs[7] [25];   // regs.v(45)
    assign n1900 = write[0] ? n876 : \regs[7] [24];   // regs.v(45)
    assign n1901 = write[0] ? n877 : \regs[7] [23];   // regs.v(45)
    assign n1902 = write[0] ? n878 : \regs[7] [22];   // regs.v(45)
    assign n1903 = write[0] ? n879 : \regs[7] [21];   // regs.v(45)
    assign n1904 = write[0] ? n880 : \regs[7] [20];   // regs.v(45)
    assign n1905 = write[0] ? n881 : \regs[7] [19];   // regs.v(45)
    assign n1906 = write[0] ? n882 : \regs[7] [18];   // regs.v(45)
    assign n1907 = write[0] ? n883 : \regs[7] [17];   // regs.v(45)
    assign n1908 = write[0] ? n884 : \regs[7] [16];   // regs.v(45)
    assign n1909 = write[0] ? n885 : \regs[7] [15];   // regs.v(45)
    assign n1910 = write[0] ? n886 : \regs[7] [14];   // regs.v(45)
    assign n1911 = write[0] ? n887 : \regs[7] [13];   // regs.v(45)
    assign n1912 = write[0] ? n888 : \regs[7] [12];   // regs.v(45)
    assign n1913 = write[0] ? n889 : \regs[7] [11];   // regs.v(45)
    assign n1914 = write[0] ? n890 : \regs[7] [10];   // regs.v(45)
    assign n1915 = write[0] ? n891 : \regs[7] [9];   // regs.v(45)
    assign n1916 = write[0] ? n892 : \regs[7] [8];   // regs.v(45)
    assign n1917 = write[0] ? n893 : \regs[7] [7];   // regs.v(45)
    assign n1918 = write[0] ? n894 : \regs[7] [6];   // regs.v(45)
    assign n1919 = write[0] ? n895 : \regs[7] [5];   // regs.v(45)
    assign n1920 = write[0] ? n896 : \regs[7] [4];   // regs.v(45)
    assign n1921 = write[0] ? n897 : \regs[7] [3];   // regs.v(45)
    assign n1922 = write[0] ? n898 : \regs[7] [2];   // regs.v(45)
    assign n1923 = write[0] ? n899 : \regs[7] [1];   // regs.v(45)
    assign n1924 = write[0] ? n900 : \regs[7] [0];   // regs.v(45)
    assign n1925 = write[0] ? n901 : \regs[6] [31];   // regs.v(45)
    assign n1926 = write[0] ? n902 : \regs[6] [30];   // regs.v(45)
    assign n1927 = write[0] ? n903 : \regs[6] [29];   // regs.v(45)
    assign n1928 = write[0] ? n904 : \regs[6] [28];   // regs.v(45)
    assign n1929 = write[0] ? n905 : \regs[6] [27];   // regs.v(45)
    assign n1930 = write[0] ? n906 : \regs[6] [26];   // regs.v(45)
    assign n1931 = write[0] ? n907 : \regs[6] [25];   // regs.v(45)
    assign n1932 = write[0] ? n908 : \regs[6] [24];   // regs.v(45)
    assign n1933 = write[0] ? n909 : \regs[6] [23];   // regs.v(45)
    assign n1934 = write[0] ? n910 : \regs[6] [22];   // regs.v(45)
    assign n1935 = write[0] ? n911 : \regs[6] [21];   // regs.v(45)
    assign n1936 = write[0] ? n912 : \regs[6] [20];   // regs.v(45)
    assign n1937 = write[0] ? n913 : \regs[6] [19];   // regs.v(45)
    assign n1938 = write[0] ? n914 : \regs[6] [18];   // regs.v(45)
    assign n1939 = write[0] ? n915 : \regs[6] [17];   // regs.v(45)
    assign n1940 = write[0] ? n916 : \regs[6] [16];   // regs.v(45)
    assign n1941 = write[0] ? n917 : \regs[6] [15];   // regs.v(45)
    assign n1942 = write[0] ? n918 : \regs[6] [14];   // regs.v(45)
    assign n1943 = write[0] ? n919 : \regs[6] [13];   // regs.v(45)
    assign n1944 = write[0] ? n920 : \regs[6] [12];   // regs.v(45)
    assign n1945 = write[0] ? n921 : \regs[6] [11];   // regs.v(45)
    assign n1946 = write[0] ? n922 : \regs[6] [10];   // regs.v(45)
    assign n1947 = write[0] ? n923 : \regs[6] [9];   // regs.v(45)
    assign n1948 = write[0] ? n924 : \regs[6] [8];   // regs.v(45)
    assign n1949 = write[0] ? n925 : \regs[6] [7];   // regs.v(45)
    assign n1950 = write[0] ? n926 : \regs[6] [6];   // regs.v(45)
    assign n1951 = write[0] ? n927 : \regs[6] [5];   // regs.v(45)
    assign n1952 = write[0] ? n928 : \regs[6] [4];   // regs.v(45)
    assign n1953 = write[0] ? n929 : \regs[6] [3];   // regs.v(45)
    assign n1954 = write[0] ? n930 : \regs[6] [2];   // regs.v(45)
    assign n1955 = write[0] ? n931 : \regs[6] [1];   // regs.v(45)
    assign n1956 = write[0] ? n932 : \regs[6] [0];   // regs.v(45)
    assign n1957 = write[0] ? n933 : \regs[5] [31];   // regs.v(45)
    assign n1958 = write[0] ? n934 : \regs[5] [30];   // regs.v(45)
    assign n1959 = write[0] ? n935 : \regs[5] [29];   // regs.v(45)
    assign n1960 = write[0] ? n936 : \regs[5] [28];   // regs.v(45)
    assign n1961 = write[0] ? n937 : \regs[5] [27];   // regs.v(45)
    assign n1962 = write[0] ? n938 : \regs[5] [26];   // regs.v(45)
    assign n1963 = write[0] ? n939 : \regs[5] [25];   // regs.v(45)
    assign n1964 = write[0] ? n940 : \regs[5] [24];   // regs.v(45)
    assign n1965 = write[0] ? n941 : \regs[5] [23];   // regs.v(45)
    assign n1966 = write[0] ? n942 : \regs[5] [22];   // regs.v(45)
    assign n1967 = write[0] ? n943 : \regs[5] [21];   // regs.v(45)
    assign n1968 = write[0] ? n944 : \regs[5] [20];   // regs.v(45)
    assign n1969 = write[0] ? n945 : \regs[5] [19];   // regs.v(45)
    assign n1970 = write[0] ? n946 : \regs[5] [18];   // regs.v(45)
    assign n1971 = write[0] ? n947 : \regs[5] [17];   // regs.v(45)
    assign n1972 = write[0] ? n948 : \regs[5] [16];   // regs.v(45)
    assign n1973 = write[0] ? n949 : \regs[5] [15];   // regs.v(45)
    assign n1974 = write[0] ? n950 : \regs[5] [14];   // regs.v(45)
    assign n1975 = write[0] ? n951 : \regs[5] [13];   // regs.v(45)
    assign n1976 = write[0] ? n952 : \regs[5] [12];   // regs.v(45)
    assign n1977 = write[0] ? n953 : \regs[5] [11];   // regs.v(45)
    assign n1978 = write[0] ? n954 : \regs[5] [10];   // regs.v(45)
    assign n1979 = write[0] ? n955 : \regs[5] [9];   // regs.v(45)
    assign n1980 = write[0] ? n956 : \regs[5] [8];   // regs.v(45)
    assign n1981 = write[0] ? n957 : \regs[5] [7];   // regs.v(45)
    assign n1982 = write[0] ? n958 : \regs[5] [6];   // regs.v(45)
    assign n1983 = write[0] ? n959 : \regs[5] [5];   // regs.v(45)
    assign n1984 = write[0] ? n960 : \regs[5] [4];   // regs.v(45)
    assign n1985 = write[0] ? n961 : \regs[5] [3];   // regs.v(45)
    assign n1986 = write[0] ? n962 : \regs[5] [2];   // regs.v(45)
    assign n1987 = write[0] ? n963 : \regs[5] [1];   // regs.v(45)
    assign n1988 = write[0] ? n964 : \regs[5] [0];   // regs.v(45)
    assign n1989 = write[0] ? n965 : \regs[4] [31];   // regs.v(45)
    assign n1990 = write[0] ? n966 : \regs[4] [30];   // regs.v(45)
    assign n1991 = write[0] ? n967 : \regs[4] [29];   // regs.v(45)
    assign n1992 = write[0] ? n968 : \regs[4] [28];   // regs.v(45)
    assign n1993 = write[0] ? n969 : \regs[4] [27];   // regs.v(45)
    assign n1994 = write[0] ? n970 : \regs[4] [26];   // regs.v(45)
    assign n1995 = write[0] ? n971 : \regs[4] [25];   // regs.v(45)
    assign n1996 = write[0] ? n972 : \regs[4] [24];   // regs.v(45)
    assign n1997 = write[0] ? n973 : \regs[4] [23];   // regs.v(45)
    assign n1998 = write[0] ? n974 : \regs[4] [22];   // regs.v(45)
    assign n1999 = write[0] ? n975 : \regs[4] [21];   // regs.v(45)
    assign n2000 = write[0] ? n976 : \regs[4] [20];   // regs.v(45)
    assign n2001 = write[0] ? n977 : \regs[4] [19];   // regs.v(45)
    assign n2002 = write[0] ? n978 : \regs[4] [18];   // regs.v(45)
    assign n2003 = write[0] ? n979 : \regs[4] [17];   // regs.v(45)
    assign n2004 = write[0] ? n980 : \regs[4] [16];   // regs.v(45)
    assign n2005 = write[0] ? n981 : \regs[4] [15];   // regs.v(45)
    assign n2006 = write[0] ? n982 : \regs[4] [14];   // regs.v(45)
    assign n2007 = write[0] ? n983 : \regs[4] [13];   // regs.v(45)
    assign n2008 = write[0] ? n984 : \regs[4] [12];   // regs.v(45)
    assign n2009 = write[0] ? n985 : \regs[4] [11];   // regs.v(45)
    assign n2010 = write[0] ? n986 : \regs[4] [10];   // regs.v(45)
    assign n2011 = write[0] ? n987 : \regs[4] [9];   // regs.v(45)
    assign n2012 = write[0] ? n988 : \regs[4] [8];   // regs.v(45)
    assign n2013 = write[0] ? n989 : \regs[4] [7];   // regs.v(45)
    assign n2014 = write[0] ? n990 : \regs[4] [6];   // regs.v(45)
    assign n2015 = write[0] ? n991 : \regs[4] [5];   // regs.v(45)
    assign n2016 = write[0] ? n992 : \regs[4] [4];   // regs.v(45)
    assign n2017 = write[0] ? n993 : \regs[4] [3];   // regs.v(45)
    assign n2018 = write[0] ? n994 : \regs[4] [2];   // regs.v(45)
    assign n2019 = write[0] ? n995 : \regs[4] [1];   // regs.v(45)
    assign n2020 = write[0] ? n996 : \regs[4] [0];   // regs.v(45)
    assign n2021 = write[0] ? n997 : \regs[3] [31];   // regs.v(45)
    assign n2022 = write[0] ? n998 : \regs[3] [30];   // regs.v(45)
    assign n2023 = write[0] ? n999 : \regs[3] [29];   // regs.v(45)
    assign n2024 = write[0] ? n1000 : \regs[3] [28];   // regs.v(45)
    assign n2025 = write[0] ? n1001 : \regs[3] [27];   // regs.v(45)
    assign n2026 = write[0] ? n1002 : \regs[3] [26];   // regs.v(45)
    assign n2027 = write[0] ? n1003 : \regs[3] [25];   // regs.v(45)
    assign n2028 = write[0] ? n1004 : \regs[3] [24];   // regs.v(45)
    assign n2029 = write[0] ? n1005 : \regs[3] [23];   // regs.v(45)
    assign n2030 = write[0] ? n1006 : \regs[3] [22];   // regs.v(45)
    assign n2031 = write[0] ? n1007 : \regs[3] [21];   // regs.v(45)
    assign n2032 = write[0] ? n1008 : \regs[3] [20];   // regs.v(45)
    assign n2033 = write[0] ? n1009 : \regs[3] [19];   // regs.v(45)
    assign n2034 = write[0] ? n1010 : \regs[3] [18];   // regs.v(45)
    assign n2035 = write[0] ? n1011 : \regs[3] [17];   // regs.v(45)
    assign n2036 = write[0] ? n1012 : \regs[3] [16];   // regs.v(45)
    assign n2037 = write[0] ? n1013 : \regs[3] [15];   // regs.v(45)
    assign n2038 = write[0] ? n1014 : \regs[3] [14];   // regs.v(45)
    assign n2039 = write[0] ? n1015 : \regs[3] [13];   // regs.v(45)
    assign n2040 = write[0] ? n1016 : \regs[3] [12];   // regs.v(45)
    assign n2041 = write[0] ? n1017 : \regs[3] [11];   // regs.v(45)
    assign n2042 = write[0] ? n1018 : \regs[3] [10];   // regs.v(45)
    assign n2043 = write[0] ? n1019 : \regs[3] [9];   // regs.v(45)
    assign n2044 = write[0] ? n1020 : \regs[3] [8];   // regs.v(45)
    assign n2045 = write[0] ? n1021 : \regs[3] [7];   // regs.v(45)
    assign n2046 = write[0] ? n1022 : \regs[3] [6];   // regs.v(45)
    assign n2047 = write[0] ? n1023 : \regs[3] [5];   // regs.v(45)
    assign n2048 = write[0] ? n1024 : \regs[3] [4];   // regs.v(45)
    assign n2049 = write[0] ? n1025 : \regs[3] [3];   // regs.v(45)
    assign n2050 = write[0] ? n1026 : \regs[3] [2];   // regs.v(45)
    assign n2051 = write[0] ? n1027 : \regs[3] [1];   // regs.v(45)
    assign n2052 = write[0] ? n1028 : \regs[3] [0];   // regs.v(45)
    assign n2053 = write[0] ? n1029 : \regs[2] [31];   // regs.v(45)
    assign n2054 = write[0] ? n1030 : \regs[2] [30];   // regs.v(45)
    assign n2055 = write[0] ? n1031 : \regs[2] [29];   // regs.v(45)
    assign n2056 = write[0] ? n1032 : \regs[2] [28];   // regs.v(45)
    assign n2057 = write[0] ? n1033 : \regs[2] [27];   // regs.v(45)
    assign n2058 = write[0] ? n1034 : \regs[2] [26];   // regs.v(45)
    assign n2059 = write[0] ? n1035 : \regs[2] [25];   // regs.v(45)
    assign n2060 = write[0] ? n1036 : \regs[2] [24];   // regs.v(45)
    assign n2061 = write[0] ? n1037 : \regs[2] [23];   // regs.v(45)
    assign n2062 = write[0] ? n1038 : \regs[2] [22];   // regs.v(45)
    assign n2063 = write[0] ? n1039 : \regs[2] [21];   // regs.v(45)
    assign n2064 = write[0] ? n1040 : \regs[2] [20];   // regs.v(45)
    assign n2065 = write[0] ? n1041 : \regs[2] [19];   // regs.v(45)
    assign n2066 = write[0] ? n1042 : \regs[2] [18];   // regs.v(45)
    assign n2067 = write[0] ? n1043 : \regs[2] [17];   // regs.v(45)
    assign n2068 = write[0] ? n1044 : \regs[2] [16];   // regs.v(45)
    assign n2069 = write[0] ? n1045 : \regs[2] [15];   // regs.v(45)
    assign n2070 = write[0] ? n1046 : \regs[2] [14];   // regs.v(45)
    assign n2071 = write[0] ? n1047 : \regs[2] [13];   // regs.v(45)
    assign n2072 = write[0] ? n1048 : \regs[2] [12];   // regs.v(45)
    assign n2073 = write[0] ? n1049 : \regs[2] [11];   // regs.v(45)
    assign n2074 = write[0] ? n1050 : \regs[2] [10];   // regs.v(45)
    assign n2075 = write[0] ? n1051 : \regs[2] [9];   // regs.v(45)
    assign n2076 = write[0] ? n1052 : \regs[2] [8];   // regs.v(45)
    assign n2077 = write[0] ? n1053 : \regs[2] [7];   // regs.v(45)
    assign n2078 = write[0] ? n1054 : \regs[2] [6];   // regs.v(45)
    assign n2079 = write[0] ? n1055 : \regs[2] [5];   // regs.v(45)
    assign n2080 = write[0] ? n1056 : \regs[2] [4];   // regs.v(45)
    assign n2081 = write[0] ? n1057 : \regs[2] [3];   // regs.v(45)
    assign n2082 = write[0] ? n1058 : \regs[2] [2];   // regs.v(45)
    assign n2083 = write[0] ? n1059 : \regs[2] [1];   // regs.v(45)
    assign n2084 = write[0] ? n1060 : \regs[2] [0];   // regs.v(45)
    assign n2085 = write[0] ? n1061 : \regs[1] [31];   // regs.v(45)
    assign n2086 = write[0] ? n1062 : \regs[1] [30];   // regs.v(45)
    assign n2087 = write[0] ? n1063 : \regs[1] [29];   // regs.v(45)
    assign n2088 = write[0] ? n1064 : \regs[1] [28];   // regs.v(45)
    assign n2089 = write[0] ? n1065 : \regs[1] [27];   // regs.v(45)
    assign n2090 = write[0] ? n1066 : \regs[1] [26];   // regs.v(45)
    assign n2091 = write[0] ? n1067 : \regs[1] [25];   // regs.v(45)
    assign n2092 = write[0] ? n1068 : \regs[1] [24];   // regs.v(45)
    assign n2093 = write[0] ? n1069 : \regs[1] [23];   // regs.v(45)
    assign n2094 = write[0] ? n1070 : \regs[1] [22];   // regs.v(45)
    assign n2095 = write[0] ? n1071 : \regs[1] [21];   // regs.v(45)
    assign n2096 = write[0] ? n1072 : \regs[1] [20];   // regs.v(45)
    assign n2097 = write[0] ? n1073 : \regs[1] [19];   // regs.v(45)
    assign n2098 = write[0] ? n1074 : \regs[1] [18];   // regs.v(45)
    assign n2099 = write[0] ? n1075 : \regs[1] [17];   // regs.v(45)
    assign n2100 = write[0] ? n1076 : \regs[1] [16];   // regs.v(45)
    assign n2101 = write[0] ? n1077 : \regs[1] [15];   // regs.v(45)
    assign n2102 = write[0] ? n1078 : \regs[1] [14];   // regs.v(45)
    assign n2103 = write[0] ? n1079 : \regs[1] [13];   // regs.v(45)
    assign n2104 = write[0] ? n1080 : \regs[1] [12];   // regs.v(45)
    assign n2105 = write[0] ? n1081 : \regs[1] [11];   // regs.v(45)
    assign n2106 = write[0] ? n1082 : \regs[1] [10];   // regs.v(45)
    assign n2107 = write[0] ? n1083 : \regs[1] [9];   // regs.v(45)
    assign n2108 = write[0] ? n1084 : \regs[1] [8];   // regs.v(45)
    assign n2109 = write[0] ? n1085 : \regs[1] [7];   // regs.v(45)
    assign n2110 = write[0] ? n1086 : \regs[1] [6];   // regs.v(45)
    assign n2111 = write[0] ? n1087 : \regs[1] [5];   // regs.v(45)
    assign n2112 = write[0] ? n1088 : \regs[1] [4];   // regs.v(45)
    assign n2113 = write[0] ? n1089 : \regs[1] [3];   // regs.v(45)
    assign n2114 = write[0] ? n1090 : \regs[1] [2];   // regs.v(45)
    assign n2115 = write[0] ? n1091 : \regs[1] [1];   // regs.v(45)
    assign n2116 = write[0] ? n1092 : \regs[1] [0];   // regs.v(45)
    assign n2117 = write[0] ? n1093 : \regs[0] [31];   // regs.v(45)
    assign n2118 = write[0] ? n1094 : \regs[0] [30];   // regs.v(45)
    assign n2119 = write[0] ? n1095 : \regs[0] [29];   // regs.v(45)
    assign n2120 = write[0] ? n1096 : \regs[0] [28];   // regs.v(45)
    assign n2121 = write[0] ? n1097 : \regs[0] [27];   // regs.v(45)
    assign n2122 = write[0] ? n1098 : \regs[0] [26];   // regs.v(45)
    assign n2123 = write[0] ? n1099 : \regs[0] [25];   // regs.v(45)
    assign n2124 = write[0] ? n1100 : \regs[0] [24];   // regs.v(45)
    assign n2125 = write[0] ? n1101 : \regs[0] [23];   // regs.v(45)
    assign n2126 = write[0] ? n1102 : \regs[0] [22];   // regs.v(45)
    assign n2127 = write[0] ? n1103 : \regs[0] [21];   // regs.v(45)
    assign n2128 = write[0] ? n1104 : \regs[0] [20];   // regs.v(45)
    assign n2129 = write[0] ? n1105 : \regs[0] [19];   // regs.v(45)
    assign n2130 = write[0] ? n1106 : \regs[0] [18];   // regs.v(45)
    assign n2131 = write[0] ? n1107 : \regs[0] [17];   // regs.v(45)
    assign n2132 = write[0] ? n1108 : \regs[0] [16];   // regs.v(45)
    assign n2133 = write[0] ? n1109 : \regs[0] [15];   // regs.v(45)
    assign n2134 = write[0] ? n1110 : \regs[0] [14];   // regs.v(45)
    assign n2135 = write[0] ? n1111 : \regs[0] [13];   // regs.v(45)
    assign n2136 = write[0] ? n1112 : \regs[0] [12];   // regs.v(45)
    assign n2137 = write[0] ? n1113 : \regs[0] [11];   // regs.v(45)
    assign n2138 = write[0] ? n1114 : \regs[0] [10];   // regs.v(45)
    assign n2139 = write[0] ? n1115 : \regs[0] [9];   // regs.v(45)
    assign n2140 = write[0] ? n1116 : \regs[0] [8];   // regs.v(45)
    assign n2141 = write[0] ? n1117 : \regs[0] [7];   // regs.v(45)
    assign n2142 = write[0] ? n1118 : \regs[0] [6];   // regs.v(45)
    assign n2143 = write[0] ? n1119 : \regs[0] [5];   // regs.v(45)
    assign n2144 = write[0] ? n1120 : \regs[0] [4];   // regs.v(45)
    assign n2145 = write[0] ? n1121 : \regs[0] [3];   // regs.v(45)
    assign n2146 = write[0] ? n1122 : \regs[0] [2];   // regs.v(45)
    assign n2147 = write[0] ? n1123 : \regs[0] [1];   // regs.v(45)
    assign n2148 = write[0] ? n1124 : \regs[0] [0];   // regs.v(45)
    Decoder_5 Decoder_2117 (.i({wa1}), .o({n2149, n2150, n2151, n2152, 
            n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, 
            n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, 
            n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, 
            n2177, n2178, n2179, n2180}));   // regs.v(46)
    assign n2181 = n2149 ? wd1[31] : n1125;   // regs.v(46)
    assign n2182 = n2149 ? wd1[30] : n1126;   // regs.v(46)
    assign n2183 = n2149 ? wd1[29] : n1127;   // regs.v(46)
    assign n2184 = n2149 ? wd1[28] : n1128;   // regs.v(46)
    assign n2185 = n2149 ? wd1[27] : n1129;   // regs.v(46)
    assign n2186 = n2149 ? wd1[26] : n1130;   // regs.v(46)
    assign n2187 = n2149 ? wd1[25] : n1131;   // regs.v(46)
    assign n2188 = n2149 ? wd1[24] : n1132;   // regs.v(46)
    assign n2189 = n2149 ? wd1[23] : n1133;   // regs.v(46)
    assign n2190 = n2149 ? wd1[22] : n1134;   // regs.v(46)
    assign n2191 = n2149 ? wd1[21] : n1135;   // regs.v(46)
    assign n2192 = n2149 ? wd1[20] : n1136;   // regs.v(46)
    assign n2193 = n2149 ? wd1[19] : n1137;   // regs.v(46)
    assign n2194 = n2149 ? wd1[18] : n1138;   // regs.v(46)
    assign n2195 = n2149 ? wd1[17] : n1139;   // regs.v(46)
    assign n2196 = n2149 ? wd1[16] : n1140;   // regs.v(46)
    assign n2197 = n2149 ? wd1[15] : n1141;   // regs.v(46)
    assign n2198 = n2149 ? wd1[14] : n1142;   // regs.v(46)
    assign n2199 = n2149 ? wd1[13] : n1143;   // regs.v(46)
    assign n2200 = n2149 ? wd1[12] : n1144;   // regs.v(46)
    assign n2201 = n2149 ? wd1[11] : n1145;   // regs.v(46)
    assign n2202 = n2149 ? wd1[10] : n1146;   // regs.v(46)
    assign n2203 = n2149 ? wd1[9] : n1147;   // regs.v(46)
    assign n2204 = n2149 ? wd1[8] : n1148;   // regs.v(46)
    assign n2205 = n2149 ? wd1[7] : n1149;   // regs.v(46)
    assign n2206 = n2149 ? wd1[6] : n1150;   // regs.v(46)
    assign n2207 = n2149 ? wd1[5] : n1151;   // regs.v(46)
    assign n2208 = n2149 ? wd1[4] : n1152;   // regs.v(46)
    assign n2209 = n2149 ? wd1[3] : n1153;   // regs.v(46)
    assign n2210 = n2149 ? wd1[2] : n1154;   // regs.v(46)
    assign n2211 = n2149 ? wd1[1] : n1155;   // regs.v(46)
    assign n2212 = n2149 ? wd1[0] : n1156;   // regs.v(46)
    assign n2213 = n2150 ? wd1[31] : n1157;   // regs.v(46)
    assign n2214 = n2150 ? wd1[30] : n1158;   // regs.v(46)
    assign n2215 = n2150 ? wd1[29] : n1159;   // regs.v(46)
    assign n2216 = n2150 ? wd1[28] : n1160;   // regs.v(46)
    assign n2217 = n2150 ? wd1[27] : n1161;   // regs.v(46)
    assign n2218 = n2150 ? wd1[26] : n1162;   // regs.v(46)
    assign n2219 = n2150 ? wd1[25] : n1163;   // regs.v(46)
    assign n2220 = n2150 ? wd1[24] : n1164;   // regs.v(46)
    assign n2221 = n2150 ? wd1[23] : n1165;   // regs.v(46)
    assign n2222 = n2150 ? wd1[22] : n1166;   // regs.v(46)
    assign n2223 = n2150 ? wd1[21] : n1167;   // regs.v(46)
    assign n2224 = n2150 ? wd1[20] : n1168;   // regs.v(46)
    assign n2225 = n2150 ? wd1[19] : n1169;   // regs.v(46)
    assign n2226 = n2150 ? wd1[18] : n1170;   // regs.v(46)
    assign n2227 = n2150 ? wd1[17] : n1171;   // regs.v(46)
    assign n2228 = n2150 ? wd1[16] : n1172;   // regs.v(46)
    assign n2229 = n2150 ? wd1[15] : n1173;   // regs.v(46)
    assign n2230 = n2150 ? wd1[14] : n1174;   // regs.v(46)
    assign n2231 = n2150 ? wd1[13] : n1175;   // regs.v(46)
    assign n2232 = n2150 ? wd1[12] : n1176;   // regs.v(46)
    assign n2233 = n2150 ? wd1[11] : n1177;   // regs.v(46)
    assign n2234 = n2150 ? wd1[10] : n1178;   // regs.v(46)
    assign n2235 = n2150 ? wd1[9] : n1179;   // regs.v(46)
    assign n2236 = n2150 ? wd1[8] : n1180;   // regs.v(46)
    assign n2237 = n2150 ? wd1[7] : n1181;   // regs.v(46)
    assign n2238 = n2150 ? wd1[6] : n1182;   // regs.v(46)
    assign n2239 = n2150 ? wd1[5] : n1183;   // regs.v(46)
    assign n2240 = n2150 ? wd1[4] : n1184;   // regs.v(46)
    assign n2241 = n2150 ? wd1[3] : n1185;   // regs.v(46)
    assign n2242 = n2150 ? wd1[2] : n1186;   // regs.v(46)
    assign n2243 = n2150 ? wd1[1] : n1187;   // regs.v(46)
    assign n2244 = n2150 ? wd1[0] : n1188;   // regs.v(46)
    assign n2245 = n2151 ? wd1[31] : n1189;   // regs.v(46)
    assign n2246 = n2151 ? wd1[30] : n1190;   // regs.v(46)
    assign n2247 = n2151 ? wd1[29] : n1191;   // regs.v(46)
    assign n2248 = n2151 ? wd1[28] : n1192;   // regs.v(46)
    assign n2249 = n2151 ? wd1[27] : n1193;   // regs.v(46)
    assign n2250 = n2151 ? wd1[26] : n1194;   // regs.v(46)
    assign n2251 = n2151 ? wd1[25] : n1195;   // regs.v(46)
    assign n2252 = n2151 ? wd1[24] : n1196;   // regs.v(46)
    assign n2253 = n2151 ? wd1[23] : n1197;   // regs.v(46)
    assign n2254 = n2151 ? wd1[22] : n1198;   // regs.v(46)
    assign n2255 = n2151 ? wd1[21] : n1199;   // regs.v(46)
    assign n2256 = n2151 ? wd1[20] : n1200;   // regs.v(46)
    assign n2257 = n2151 ? wd1[19] : n1201;   // regs.v(46)
    assign n2258 = n2151 ? wd1[18] : n1202;   // regs.v(46)
    assign n2259 = n2151 ? wd1[17] : n1203;   // regs.v(46)
    assign n2260 = n2151 ? wd1[16] : n1204;   // regs.v(46)
    assign n2261 = n2151 ? wd1[15] : n1205;   // regs.v(46)
    assign n2262 = n2151 ? wd1[14] : n1206;   // regs.v(46)
    assign n2263 = n2151 ? wd1[13] : n1207;   // regs.v(46)
    assign n2264 = n2151 ? wd1[12] : n1208;   // regs.v(46)
    assign n2265 = n2151 ? wd1[11] : n1209;   // regs.v(46)
    assign n2266 = n2151 ? wd1[10] : n1210;   // regs.v(46)
    assign n2267 = n2151 ? wd1[9] : n1211;   // regs.v(46)
    assign n2268 = n2151 ? wd1[8] : n1212;   // regs.v(46)
    assign n2269 = n2151 ? wd1[7] : n1213;   // regs.v(46)
    assign n2270 = n2151 ? wd1[6] : n1214;   // regs.v(46)
    assign n2271 = n2151 ? wd1[5] : n1215;   // regs.v(46)
    assign n2272 = n2151 ? wd1[4] : n1216;   // regs.v(46)
    assign n2273 = n2151 ? wd1[3] : n1217;   // regs.v(46)
    assign n2274 = n2151 ? wd1[2] : n1218;   // regs.v(46)
    assign n2275 = n2151 ? wd1[1] : n1219;   // regs.v(46)
    assign n2276 = n2151 ? wd1[0] : n1220;   // regs.v(46)
    assign n2277 = n2152 ? wd1[31] : n1221;   // regs.v(46)
    assign n2278 = n2152 ? wd1[30] : n1222;   // regs.v(46)
    assign n2279 = n2152 ? wd1[29] : n1223;   // regs.v(46)
    assign n2280 = n2152 ? wd1[28] : n1224;   // regs.v(46)
    assign n2281 = n2152 ? wd1[27] : n1225;   // regs.v(46)
    assign n2282 = n2152 ? wd1[26] : n1226;   // regs.v(46)
    assign n2283 = n2152 ? wd1[25] : n1227;   // regs.v(46)
    assign n2284 = n2152 ? wd1[24] : n1228;   // regs.v(46)
    assign n2285 = n2152 ? wd1[23] : n1229;   // regs.v(46)
    assign n2286 = n2152 ? wd1[22] : n1230;   // regs.v(46)
    assign n2287 = n2152 ? wd1[21] : n1231;   // regs.v(46)
    assign n2288 = n2152 ? wd1[20] : n1232;   // regs.v(46)
    assign n2289 = n2152 ? wd1[19] : n1233;   // regs.v(46)
    assign n2290 = n2152 ? wd1[18] : n1234;   // regs.v(46)
    assign n2291 = n2152 ? wd1[17] : n1235;   // regs.v(46)
    assign n2292 = n2152 ? wd1[16] : n1236;   // regs.v(46)
    assign n2293 = n2152 ? wd1[15] : n1237;   // regs.v(46)
    assign n2294 = n2152 ? wd1[14] : n1238;   // regs.v(46)
    assign n2295 = n2152 ? wd1[13] : n1239;   // regs.v(46)
    assign n2296 = n2152 ? wd1[12] : n1240;   // regs.v(46)
    assign n2297 = n2152 ? wd1[11] : n1241;   // regs.v(46)
    assign n2298 = n2152 ? wd1[10] : n1242;   // regs.v(46)
    assign n2299 = n2152 ? wd1[9] : n1243;   // regs.v(46)
    assign n2300 = n2152 ? wd1[8] : n1244;   // regs.v(46)
    assign n2301 = n2152 ? wd1[7] : n1245;   // regs.v(46)
    assign n2302 = n2152 ? wd1[6] : n1246;   // regs.v(46)
    assign n2303 = n2152 ? wd1[5] : n1247;   // regs.v(46)
    assign n2304 = n2152 ? wd1[4] : n1248;   // regs.v(46)
    assign n2305 = n2152 ? wd1[3] : n1249;   // regs.v(46)
    assign n2306 = n2152 ? wd1[2] : n1250;   // regs.v(46)
    assign n2307 = n2152 ? wd1[1] : n1251;   // regs.v(46)
    assign n2308 = n2152 ? wd1[0] : n1252;   // regs.v(46)
    assign n2309 = n2153 ? wd1[31] : n1253;   // regs.v(46)
    assign n2310 = n2153 ? wd1[30] : n1254;   // regs.v(46)
    assign n2311 = n2153 ? wd1[29] : n1255;   // regs.v(46)
    assign n2312 = n2153 ? wd1[28] : n1256;   // regs.v(46)
    assign n2313 = n2153 ? wd1[27] : n1257;   // regs.v(46)
    assign n2314 = n2153 ? wd1[26] : n1258;   // regs.v(46)
    assign n2315 = n2153 ? wd1[25] : n1259;   // regs.v(46)
    assign n2316 = n2153 ? wd1[24] : n1260;   // regs.v(46)
    assign n2317 = n2153 ? wd1[23] : n1261;   // regs.v(46)
    assign n2318 = n2153 ? wd1[22] : n1262;   // regs.v(46)
    assign n2319 = n2153 ? wd1[21] : n1263;   // regs.v(46)
    assign n2320 = n2153 ? wd1[20] : n1264;   // regs.v(46)
    assign n2321 = n2153 ? wd1[19] : n1265;   // regs.v(46)
    assign n2322 = n2153 ? wd1[18] : n1266;   // regs.v(46)
    assign n2323 = n2153 ? wd1[17] : n1267;   // regs.v(46)
    assign n2324 = n2153 ? wd1[16] : n1268;   // regs.v(46)
    assign n2325 = n2153 ? wd1[15] : n1269;   // regs.v(46)
    assign n2326 = n2153 ? wd1[14] : n1270;   // regs.v(46)
    assign n2327 = n2153 ? wd1[13] : n1271;   // regs.v(46)
    assign n2328 = n2153 ? wd1[12] : n1272;   // regs.v(46)
    assign n2329 = n2153 ? wd1[11] : n1273;   // regs.v(46)
    assign n2330 = n2153 ? wd1[10] : n1274;   // regs.v(46)
    assign n2331 = n2153 ? wd1[9] : n1275;   // regs.v(46)
    assign n2332 = n2153 ? wd1[8] : n1276;   // regs.v(46)
    assign n2333 = n2153 ? wd1[7] : n1277;   // regs.v(46)
    assign n2334 = n2153 ? wd1[6] : n1278;   // regs.v(46)
    assign n2335 = n2153 ? wd1[5] : n1279;   // regs.v(46)
    assign n2336 = n2153 ? wd1[4] : n1280;   // regs.v(46)
    assign n2337 = n2153 ? wd1[3] : n1281;   // regs.v(46)
    assign n2338 = n2153 ? wd1[2] : n1282;   // regs.v(46)
    assign n2339 = n2153 ? wd1[1] : n1283;   // regs.v(46)
    assign n2340 = n2153 ? wd1[0] : n1284;   // regs.v(46)
    assign n2341 = n2154 ? wd1[31] : n1285;   // regs.v(46)
    assign n2342 = n2154 ? wd1[30] : n1286;   // regs.v(46)
    assign n2343 = n2154 ? wd1[29] : n1287;   // regs.v(46)
    assign n2344 = n2154 ? wd1[28] : n1288;   // regs.v(46)
    assign n2345 = n2154 ? wd1[27] : n1289;   // regs.v(46)
    assign n2346 = n2154 ? wd1[26] : n1290;   // regs.v(46)
    assign n2347 = n2154 ? wd1[25] : n1291;   // regs.v(46)
    assign n2348 = n2154 ? wd1[24] : n1292;   // regs.v(46)
    assign n2349 = n2154 ? wd1[23] : n1293;   // regs.v(46)
    assign n2350 = n2154 ? wd1[22] : n1294;   // regs.v(46)
    assign n2351 = n2154 ? wd1[21] : n1295;   // regs.v(46)
    assign n2352 = n2154 ? wd1[20] : n1296;   // regs.v(46)
    assign n2353 = n2154 ? wd1[19] : n1297;   // regs.v(46)
    assign n2354 = n2154 ? wd1[18] : n1298;   // regs.v(46)
    assign n2355 = n2154 ? wd1[17] : n1299;   // regs.v(46)
    assign n2356 = n2154 ? wd1[16] : n1300;   // regs.v(46)
    assign n2357 = n2154 ? wd1[15] : n1301;   // regs.v(46)
    assign n2358 = n2154 ? wd1[14] : n1302;   // regs.v(46)
    assign n2359 = n2154 ? wd1[13] : n1303;   // regs.v(46)
    assign n2360 = n2154 ? wd1[12] : n1304;   // regs.v(46)
    assign n2361 = n2154 ? wd1[11] : n1305;   // regs.v(46)
    assign n2362 = n2154 ? wd1[10] : n1306;   // regs.v(46)
    assign n2363 = n2154 ? wd1[9] : n1307;   // regs.v(46)
    assign n2364 = n2154 ? wd1[8] : n1308;   // regs.v(46)
    assign n2365 = n2154 ? wd1[7] : n1309;   // regs.v(46)
    assign n2366 = n2154 ? wd1[6] : n1310;   // regs.v(46)
    assign n2367 = n2154 ? wd1[5] : n1311;   // regs.v(46)
    assign n2368 = n2154 ? wd1[4] : n1312;   // regs.v(46)
    assign n2369 = n2154 ? wd1[3] : n1313;   // regs.v(46)
    assign n2370 = n2154 ? wd1[2] : n1314;   // regs.v(46)
    assign n2371 = n2154 ? wd1[1] : n1315;   // regs.v(46)
    assign n2372 = n2154 ? wd1[0] : n1316;   // regs.v(46)
    assign n2373 = n2155 ? wd1[31] : n1317;   // regs.v(46)
    assign n2374 = n2155 ? wd1[30] : n1318;   // regs.v(46)
    assign n2375 = n2155 ? wd1[29] : n1319;   // regs.v(46)
    assign n2376 = n2155 ? wd1[28] : n1320;   // regs.v(46)
    assign n2377 = n2155 ? wd1[27] : n1321;   // regs.v(46)
    assign n2378 = n2155 ? wd1[26] : n1322;   // regs.v(46)
    assign n2379 = n2155 ? wd1[25] : n1323;   // regs.v(46)
    assign n2380 = n2155 ? wd1[24] : n1324;   // regs.v(46)
    assign n2381 = n2155 ? wd1[23] : n1325;   // regs.v(46)
    assign n2382 = n2155 ? wd1[22] : n1326;   // regs.v(46)
    assign n2383 = n2155 ? wd1[21] : n1327;   // regs.v(46)
    assign n2384 = n2155 ? wd1[20] : n1328;   // regs.v(46)
    assign n2385 = n2155 ? wd1[19] : n1329;   // regs.v(46)
    assign n2386 = n2155 ? wd1[18] : n1330;   // regs.v(46)
    assign n2387 = n2155 ? wd1[17] : n1331;   // regs.v(46)
    assign n2388 = n2155 ? wd1[16] : n1332;   // regs.v(46)
    assign n2389 = n2155 ? wd1[15] : n1333;   // regs.v(46)
    assign n2390 = n2155 ? wd1[14] : n1334;   // regs.v(46)
    assign n2391 = n2155 ? wd1[13] : n1335;   // regs.v(46)
    assign n2392 = n2155 ? wd1[12] : n1336;   // regs.v(46)
    assign n2393 = n2155 ? wd1[11] : n1337;   // regs.v(46)
    assign n2394 = n2155 ? wd1[10] : n1338;   // regs.v(46)
    assign n2395 = n2155 ? wd1[9] : n1339;   // regs.v(46)
    assign n2396 = n2155 ? wd1[8] : n1340;   // regs.v(46)
    assign n2397 = n2155 ? wd1[7] : n1341;   // regs.v(46)
    assign n2398 = n2155 ? wd1[6] : n1342;   // regs.v(46)
    assign n2399 = n2155 ? wd1[5] : n1343;   // regs.v(46)
    assign n2400 = n2155 ? wd1[4] : n1344;   // regs.v(46)
    assign n2401 = n2155 ? wd1[3] : n1345;   // regs.v(46)
    assign n2402 = n2155 ? wd1[2] : n1346;   // regs.v(46)
    assign n2403 = n2155 ? wd1[1] : n1347;   // regs.v(46)
    assign n2404 = n2155 ? wd1[0] : n1348;   // regs.v(46)
    assign n2405 = n2156 ? wd1[31] : n1349;   // regs.v(46)
    assign n2406 = n2156 ? wd1[30] : n1350;   // regs.v(46)
    assign n2407 = n2156 ? wd1[29] : n1351;   // regs.v(46)
    assign n2408 = n2156 ? wd1[28] : n1352;   // regs.v(46)
    assign n2409 = n2156 ? wd1[27] : n1353;   // regs.v(46)
    assign n2410 = n2156 ? wd1[26] : n1354;   // regs.v(46)
    assign n2411 = n2156 ? wd1[25] : n1355;   // regs.v(46)
    assign n2412 = n2156 ? wd1[24] : n1356;   // regs.v(46)
    assign n2413 = n2156 ? wd1[23] : n1357;   // regs.v(46)
    assign n2414 = n2156 ? wd1[22] : n1358;   // regs.v(46)
    assign n2415 = n2156 ? wd1[21] : n1359;   // regs.v(46)
    assign n2416 = n2156 ? wd1[20] : n1360;   // regs.v(46)
    assign n2417 = n2156 ? wd1[19] : n1361;   // regs.v(46)
    assign n2418 = n2156 ? wd1[18] : n1362;   // regs.v(46)
    assign n2419 = n2156 ? wd1[17] : n1363;   // regs.v(46)
    assign n2420 = n2156 ? wd1[16] : n1364;   // regs.v(46)
    assign n2421 = n2156 ? wd1[15] : n1365;   // regs.v(46)
    assign n2422 = n2156 ? wd1[14] : n1366;   // regs.v(46)
    assign n2423 = n2156 ? wd1[13] : n1367;   // regs.v(46)
    assign n2424 = n2156 ? wd1[12] : n1368;   // regs.v(46)
    assign n2425 = n2156 ? wd1[11] : n1369;   // regs.v(46)
    assign n2426 = n2156 ? wd1[10] : n1370;   // regs.v(46)
    assign n2427 = n2156 ? wd1[9] : n1371;   // regs.v(46)
    assign n2428 = n2156 ? wd1[8] : n1372;   // regs.v(46)
    assign n2429 = n2156 ? wd1[7] : n1373;   // regs.v(46)
    assign n2430 = n2156 ? wd1[6] : n1374;   // regs.v(46)
    assign n2431 = n2156 ? wd1[5] : n1375;   // regs.v(46)
    assign n2432 = n2156 ? wd1[4] : n1376;   // regs.v(46)
    assign n2433 = n2156 ? wd1[3] : n1377;   // regs.v(46)
    assign n2434 = n2156 ? wd1[2] : n1378;   // regs.v(46)
    assign n2435 = n2156 ? wd1[1] : n1379;   // regs.v(46)
    assign n2436 = n2156 ? wd1[0] : n1380;   // regs.v(46)
    assign n2437 = n2157 ? wd1[31] : n1381;   // regs.v(46)
    assign n2438 = n2157 ? wd1[30] : n1382;   // regs.v(46)
    assign n2439 = n2157 ? wd1[29] : n1383;   // regs.v(46)
    assign n2440 = n2157 ? wd1[28] : n1384;   // regs.v(46)
    assign n2441 = n2157 ? wd1[27] : n1385;   // regs.v(46)
    assign n2442 = n2157 ? wd1[26] : n1386;   // regs.v(46)
    assign n2443 = n2157 ? wd1[25] : n1387;   // regs.v(46)
    assign n2444 = n2157 ? wd1[24] : n1388;   // regs.v(46)
    assign n2445 = n2157 ? wd1[23] : n1389;   // regs.v(46)
    assign n2446 = n2157 ? wd1[22] : n1390;   // regs.v(46)
    assign n2447 = n2157 ? wd1[21] : n1391;   // regs.v(46)
    assign n2448 = n2157 ? wd1[20] : n1392;   // regs.v(46)
    assign n2449 = n2157 ? wd1[19] : n1393;   // regs.v(46)
    assign n2450 = n2157 ? wd1[18] : n1394;   // regs.v(46)
    assign n2451 = n2157 ? wd1[17] : n1395;   // regs.v(46)
    assign n2452 = n2157 ? wd1[16] : n1396;   // regs.v(46)
    assign n2453 = n2157 ? wd1[15] : n1397;   // regs.v(46)
    assign n2454 = n2157 ? wd1[14] : n1398;   // regs.v(46)
    assign n2455 = n2157 ? wd1[13] : n1399;   // regs.v(46)
    assign n2456 = n2157 ? wd1[12] : n1400;   // regs.v(46)
    assign n2457 = n2157 ? wd1[11] : n1401;   // regs.v(46)
    assign n2458 = n2157 ? wd1[10] : n1402;   // regs.v(46)
    assign n2459 = n2157 ? wd1[9] : n1403;   // regs.v(46)
    assign n2460 = n2157 ? wd1[8] : n1404;   // regs.v(46)
    assign n2461 = n2157 ? wd1[7] : n1405;   // regs.v(46)
    assign n2462 = n2157 ? wd1[6] : n1406;   // regs.v(46)
    assign n2463 = n2157 ? wd1[5] : n1407;   // regs.v(46)
    assign n2464 = n2157 ? wd1[4] : n1408;   // regs.v(46)
    assign n2465 = n2157 ? wd1[3] : n1409;   // regs.v(46)
    assign n2466 = n2157 ? wd1[2] : n1410;   // regs.v(46)
    assign n2467 = n2157 ? wd1[1] : n1411;   // regs.v(46)
    assign n2468 = n2157 ? wd1[0] : n1412;   // regs.v(46)
    assign n2469 = n2158 ? wd1[31] : n1413;   // regs.v(46)
    assign n2470 = n2158 ? wd1[30] : n1414;   // regs.v(46)
    assign n2471 = n2158 ? wd1[29] : n1415;   // regs.v(46)
    assign n2472 = n2158 ? wd1[28] : n1416;   // regs.v(46)
    assign n2473 = n2158 ? wd1[27] : n1417;   // regs.v(46)
    assign n2474 = n2158 ? wd1[26] : n1418;   // regs.v(46)
    assign n2475 = n2158 ? wd1[25] : n1419;   // regs.v(46)
    assign n2476 = n2158 ? wd1[24] : n1420;   // regs.v(46)
    assign n2477 = n2158 ? wd1[23] : n1421;   // regs.v(46)
    assign n2478 = n2158 ? wd1[22] : n1422;   // regs.v(46)
    assign n2479 = n2158 ? wd1[21] : n1423;   // regs.v(46)
    assign n2480 = n2158 ? wd1[20] : n1424;   // regs.v(46)
    assign n2481 = n2158 ? wd1[19] : n1425;   // regs.v(46)
    assign n2482 = n2158 ? wd1[18] : n1426;   // regs.v(46)
    assign n2483 = n2158 ? wd1[17] : n1427;   // regs.v(46)
    assign n2484 = n2158 ? wd1[16] : n1428;   // regs.v(46)
    assign n2485 = n2158 ? wd1[15] : n1429;   // regs.v(46)
    assign n2486 = n2158 ? wd1[14] : n1430;   // regs.v(46)
    assign n2487 = n2158 ? wd1[13] : n1431;   // regs.v(46)
    assign n2488 = n2158 ? wd1[12] : n1432;   // regs.v(46)
    assign n2489 = n2158 ? wd1[11] : n1433;   // regs.v(46)
    assign n2490 = n2158 ? wd1[10] : n1434;   // regs.v(46)
    assign n2491 = n2158 ? wd1[9] : n1435;   // regs.v(46)
    assign n2492 = n2158 ? wd1[8] : n1436;   // regs.v(46)
    assign n2493 = n2158 ? wd1[7] : n1437;   // regs.v(46)
    assign n2494 = n2158 ? wd1[6] : n1438;   // regs.v(46)
    assign n2495 = n2158 ? wd1[5] : n1439;   // regs.v(46)
    assign n2496 = n2158 ? wd1[4] : n1440;   // regs.v(46)
    assign n2497 = n2158 ? wd1[3] : n1441;   // regs.v(46)
    assign n2498 = n2158 ? wd1[2] : n1442;   // regs.v(46)
    assign n2499 = n2158 ? wd1[1] : n1443;   // regs.v(46)
    assign n2500 = n2158 ? wd1[0] : n1444;   // regs.v(46)
    assign n2501 = n2159 ? wd1[31] : n1445;   // regs.v(46)
    assign n2502 = n2159 ? wd1[30] : n1446;   // regs.v(46)
    assign n2503 = n2159 ? wd1[29] : n1447;   // regs.v(46)
    assign n2504 = n2159 ? wd1[28] : n1448;   // regs.v(46)
    assign n2505 = n2159 ? wd1[27] : n1449;   // regs.v(46)
    assign n2506 = n2159 ? wd1[26] : n1450;   // regs.v(46)
    assign n2507 = n2159 ? wd1[25] : n1451;   // regs.v(46)
    assign n2508 = n2159 ? wd1[24] : n1452;   // regs.v(46)
    assign n2509 = n2159 ? wd1[23] : n1453;   // regs.v(46)
    assign n2510 = n2159 ? wd1[22] : n1454;   // regs.v(46)
    assign n2511 = n2159 ? wd1[21] : n1455;   // regs.v(46)
    assign n2512 = n2159 ? wd1[20] : n1456;   // regs.v(46)
    assign n2513 = n2159 ? wd1[19] : n1457;   // regs.v(46)
    assign n2514 = n2159 ? wd1[18] : n1458;   // regs.v(46)
    assign n2515 = n2159 ? wd1[17] : n1459;   // regs.v(46)
    assign n2516 = n2159 ? wd1[16] : n1460;   // regs.v(46)
    assign n2517 = n2159 ? wd1[15] : n1461;   // regs.v(46)
    assign n2518 = n2159 ? wd1[14] : n1462;   // regs.v(46)
    assign n2519 = n2159 ? wd1[13] : n1463;   // regs.v(46)
    assign n2520 = n2159 ? wd1[12] : n1464;   // regs.v(46)
    assign n2521 = n2159 ? wd1[11] : n1465;   // regs.v(46)
    assign n2522 = n2159 ? wd1[10] : n1466;   // regs.v(46)
    assign n2523 = n2159 ? wd1[9] : n1467;   // regs.v(46)
    assign n2524 = n2159 ? wd1[8] : n1468;   // regs.v(46)
    assign n2525 = n2159 ? wd1[7] : n1469;   // regs.v(46)
    assign n2526 = n2159 ? wd1[6] : n1470;   // regs.v(46)
    assign n2527 = n2159 ? wd1[5] : n1471;   // regs.v(46)
    assign n2528 = n2159 ? wd1[4] : n1472;   // regs.v(46)
    assign n2529 = n2159 ? wd1[3] : n1473;   // regs.v(46)
    assign n2530 = n2159 ? wd1[2] : n1474;   // regs.v(46)
    assign n2531 = n2159 ? wd1[1] : n1475;   // regs.v(46)
    assign n2532 = n2159 ? wd1[0] : n1476;   // regs.v(46)
    assign n2533 = n2160 ? wd1[31] : n1477;   // regs.v(46)
    assign n2534 = n2160 ? wd1[30] : n1478;   // regs.v(46)
    assign n2535 = n2160 ? wd1[29] : n1479;   // regs.v(46)
    assign n2536 = n2160 ? wd1[28] : n1480;   // regs.v(46)
    assign n2537 = n2160 ? wd1[27] : n1481;   // regs.v(46)
    assign n2538 = n2160 ? wd1[26] : n1482;   // regs.v(46)
    assign n2539 = n2160 ? wd1[25] : n1483;   // regs.v(46)
    assign n2540 = n2160 ? wd1[24] : n1484;   // regs.v(46)
    assign n2541 = n2160 ? wd1[23] : n1485;   // regs.v(46)
    assign n2542 = n2160 ? wd1[22] : n1486;   // regs.v(46)
    assign n2543 = n2160 ? wd1[21] : n1487;   // regs.v(46)
    assign n2544 = n2160 ? wd1[20] : n1488;   // regs.v(46)
    assign n2545 = n2160 ? wd1[19] : n1489;   // regs.v(46)
    assign n2546 = n2160 ? wd1[18] : n1490;   // regs.v(46)
    assign n2547 = n2160 ? wd1[17] : n1491;   // regs.v(46)
    assign n2548 = n2160 ? wd1[16] : n1492;   // regs.v(46)
    assign n2549 = n2160 ? wd1[15] : n1493;   // regs.v(46)
    assign n2550 = n2160 ? wd1[14] : n1494;   // regs.v(46)
    assign n2551 = n2160 ? wd1[13] : n1495;   // regs.v(46)
    assign n2552 = n2160 ? wd1[12] : n1496;   // regs.v(46)
    assign n2553 = n2160 ? wd1[11] : n1497;   // regs.v(46)
    assign n2554 = n2160 ? wd1[10] : n1498;   // regs.v(46)
    assign n2555 = n2160 ? wd1[9] : n1499;   // regs.v(46)
    assign n2556 = n2160 ? wd1[8] : n1500;   // regs.v(46)
    assign n2557 = n2160 ? wd1[7] : n1501;   // regs.v(46)
    assign n2558 = n2160 ? wd1[6] : n1502;   // regs.v(46)
    assign n2559 = n2160 ? wd1[5] : n1503;   // regs.v(46)
    assign n2560 = n2160 ? wd1[4] : n1504;   // regs.v(46)
    assign n2561 = n2160 ? wd1[3] : n1505;   // regs.v(46)
    assign n2562 = n2160 ? wd1[2] : n1506;   // regs.v(46)
    assign n2563 = n2160 ? wd1[1] : n1507;   // regs.v(46)
    assign n2564 = n2160 ? wd1[0] : n1508;   // regs.v(46)
    assign n2565 = n2161 ? wd1[31] : n1509;   // regs.v(46)
    assign n2566 = n2161 ? wd1[30] : n1510;   // regs.v(46)
    assign n2567 = n2161 ? wd1[29] : n1511;   // regs.v(46)
    assign n2568 = n2161 ? wd1[28] : n1512;   // regs.v(46)
    assign n2569 = n2161 ? wd1[27] : n1513;   // regs.v(46)
    assign n2570 = n2161 ? wd1[26] : n1514;   // regs.v(46)
    assign n2571 = n2161 ? wd1[25] : n1515;   // regs.v(46)
    assign n2572 = n2161 ? wd1[24] : n1516;   // regs.v(46)
    assign n2573 = n2161 ? wd1[23] : n1517;   // regs.v(46)
    assign n2574 = n2161 ? wd1[22] : n1518;   // regs.v(46)
    assign n2575 = n2161 ? wd1[21] : n1519;   // regs.v(46)
    assign n2576 = n2161 ? wd1[20] : n1520;   // regs.v(46)
    assign n2577 = n2161 ? wd1[19] : n1521;   // regs.v(46)
    assign n2578 = n2161 ? wd1[18] : n1522;   // regs.v(46)
    assign n2579 = n2161 ? wd1[17] : n1523;   // regs.v(46)
    assign n2580 = n2161 ? wd1[16] : n1524;   // regs.v(46)
    assign n2581 = n2161 ? wd1[15] : n1525;   // regs.v(46)
    assign n2582 = n2161 ? wd1[14] : n1526;   // regs.v(46)
    assign n2583 = n2161 ? wd1[13] : n1527;   // regs.v(46)
    assign n2584 = n2161 ? wd1[12] : n1528;   // regs.v(46)
    assign n2585 = n2161 ? wd1[11] : n1529;   // regs.v(46)
    assign n2586 = n2161 ? wd1[10] : n1530;   // regs.v(46)
    assign n2587 = n2161 ? wd1[9] : n1531;   // regs.v(46)
    assign n2588 = n2161 ? wd1[8] : n1532;   // regs.v(46)
    assign n2589 = n2161 ? wd1[7] : n1533;   // regs.v(46)
    assign n2590 = n2161 ? wd1[6] : n1534;   // regs.v(46)
    assign n2591 = n2161 ? wd1[5] : n1535;   // regs.v(46)
    assign n2592 = n2161 ? wd1[4] : n1536;   // regs.v(46)
    assign n2593 = n2161 ? wd1[3] : n1537;   // regs.v(46)
    assign n2594 = n2161 ? wd1[2] : n1538;   // regs.v(46)
    assign n2595 = n2161 ? wd1[1] : n1539;   // regs.v(46)
    assign n2596 = n2161 ? wd1[0] : n1540;   // regs.v(46)
    assign n2597 = n2162 ? wd1[31] : n1541;   // regs.v(46)
    assign n2598 = n2162 ? wd1[30] : n1542;   // regs.v(46)
    assign n2599 = n2162 ? wd1[29] : n1543;   // regs.v(46)
    assign n2600 = n2162 ? wd1[28] : n1544;   // regs.v(46)
    assign n2601 = n2162 ? wd1[27] : n1545;   // regs.v(46)
    assign n2602 = n2162 ? wd1[26] : n1546;   // regs.v(46)
    assign n2603 = n2162 ? wd1[25] : n1547;   // regs.v(46)
    assign n2604 = n2162 ? wd1[24] : n1548;   // regs.v(46)
    assign n2605 = n2162 ? wd1[23] : n1549;   // regs.v(46)
    assign n2606 = n2162 ? wd1[22] : n1550;   // regs.v(46)
    assign n2607 = n2162 ? wd1[21] : n1551;   // regs.v(46)
    assign n2608 = n2162 ? wd1[20] : n1552;   // regs.v(46)
    assign n2609 = n2162 ? wd1[19] : n1553;   // regs.v(46)
    assign n2610 = n2162 ? wd1[18] : n1554;   // regs.v(46)
    assign n2611 = n2162 ? wd1[17] : n1555;   // regs.v(46)
    assign n2612 = n2162 ? wd1[16] : n1556;   // regs.v(46)
    assign n2613 = n2162 ? wd1[15] : n1557;   // regs.v(46)
    assign n2614 = n2162 ? wd1[14] : n1558;   // regs.v(46)
    assign n2615 = n2162 ? wd1[13] : n1559;   // regs.v(46)
    assign n2616 = n2162 ? wd1[12] : n1560;   // regs.v(46)
    assign n2617 = n2162 ? wd1[11] : n1561;   // regs.v(46)
    assign n2618 = n2162 ? wd1[10] : n1562;   // regs.v(46)
    assign n2619 = n2162 ? wd1[9] : n1563;   // regs.v(46)
    assign n2620 = n2162 ? wd1[8] : n1564;   // regs.v(46)
    assign n2621 = n2162 ? wd1[7] : n1565;   // regs.v(46)
    assign n2622 = n2162 ? wd1[6] : n1566;   // regs.v(46)
    assign n2623 = n2162 ? wd1[5] : n1567;   // regs.v(46)
    assign n2624 = n2162 ? wd1[4] : n1568;   // regs.v(46)
    assign n2625 = n2162 ? wd1[3] : n1569;   // regs.v(46)
    assign n2626 = n2162 ? wd1[2] : n1570;   // regs.v(46)
    assign n2627 = n2162 ? wd1[1] : n1571;   // regs.v(46)
    assign n2628 = n2162 ? wd1[0] : n1572;   // regs.v(46)
    assign n2629 = n2163 ? wd1[31] : n1573;   // regs.v(46)
    assign n2630 = n2163 ? wd1[30] : n1574;   // regs.v(46)
    assign n2631 = n2163 ? wd1[29] : n1575;   // regs.v(46)
    assign n2632 = n2163 ? wd1[28] : n1576;   // regs.v(46)
    assign n2633 = n2163 ? wd1[27] : n1577;   // regs.v(46)
    assign n2634 = n2163 ? wd1[26] : n1578;   // regs.v(46)
    assign n2635 = n2163 ? wd1[25] : n1579;   // regs.v(46)
    assign n2636 = n2163 ? wd1[24] : n1580;   // regs.v(46)
    assign n2637 = n2163 ? wd1[23] : n1581;   // regs.v(46)
    assign n2638 = n2163 ? wd1[22] : n1582;   // regs.v(46)
    assign n2639 = n2163 ? wd1[21] : n1583;   // regs.v(46)
    assign n2640 = n2163 ? wd1[20] : n1584;   // regs.v(46)
    assign n2641 = n2163 ? wd1[19] : n1585;   // regs.v(46)
    assign n2642 = n2163 ? wd1[18] : n1586;   // regs.v(46)
    assign n2643 = n2163 ? wd1[17] : n1587;   // regs.v(46)
    assign n2644 = n2163 ? wd1[16] : n1588;   // regs.v(46)
    assign n2645 = n2163 ? wd1[15] : n1589;   // regs.v(46)
    assign n2646 = n2163 ? wd1[14] : n1590;   // regs.v(46)
    assign n2647 = n2163 ? wd1[13] : n1591;   // regs.v(46)
    assign n2648 = n2163 ? wd1[12] : n1592;   // regs.v(46)
    assign n2649 = n2163 ? wd1[11] : n1593;   // regs.v(46)
    assign n2650 = n2163 ? wd1[10] : n1594;   // regs.v(46)
    assign n2651 = n2163 ? wd1[9] : n1595;   // regs.v(46)
    assign n2652 = n2163 ? wd1[8] : n1596;   // regs.v(46)
    assign n2653 = n2163 ? wd1[7] : n1597;   // regs.v(46)
    assign n2654 = n2163 ? wd1[6] : n1598;   // regs.v(46)
    assign n2655 = n2163 ? wd1[5] : n1599;   // regs.v(46)
    assign n2656 = n2163 ? wd1[4] : n1600;   // regs.v(46)
    assign n2657 = n2163 ? wd1[3] : n1601;   // regs.v(46)
    assign n2658 = n2163 ? wd1[2] : n1602;   // regs.v(46)
    assign n2659 = n2163 ? wd1[1] : n1603;   // regs.v(46)
    assign n2660 = n2163 ? wd1[0] : n1604;   // regs.v(46)
    assign n2661 = n2164 ? wd1[31] : n1605;   // regs.v(46)
    assign n2662 = n2164 ? wd1[30] : n1606;   // regs.v(46)
    assign n2663 = n2164 ? wd1[29] : n1607;   // regs.v(46)
    assign n2664 = n2164 ? wd1[28] : n1608;   // regs.v(46)
    assign n2665 = n2164 ? wd1[27] : n1609;   // regs.v(46)
    assign n2666 = n2164 ? wd1[26] : n1610;   // regs.v(46)
    assign n2667 = n2164 ? wd1[25] : n1611;   // regs.v(46)
    assign n2668 = n2164 ? wd1[24] : n1612;   // regs.v(46)
    assign n2669 = n2164 ? wd1[23] : n1613;   // regs.v(46)
    assign n2670 = n2164 ? wd1[22] : n1614;   // regs.v(46)
    assign n2671 = n2164 ? wd1[21] : n1615;   // regs.v(46)
    assign n2672 = n2164 ? wd1[20] : n1616;   // regs.v(46)
    assign n2673 = n2164 ? wd1[19] : n1617;   // regs.v(46)
    assign n2674 = n2164 ? wd1[18] : n1618;   // regs.v(46)
    assign n2675 = n2164 ? wd1[17] : n1619;   // regs.v(46)
    assign n2676 = n2164 ? wd1[16] : n1620;   // regs.v(46)
    assign n2677 = n2164 ? wd1[15] : n1621;   // regs.v(46)
    assign n2678 = n2164 ? wd1[14] : n1622;   // regs.v(46)
    assign n2679 = n2164 ? wd1[13] : n1623;   // regs.v(46)
    assign n2680 = n2164 ? wd1[12] : n1624;   // regs.v(46)
    assign n2681 = n2164 ? wd1[11] : n1625;   // regs.v(46)
    assign n2682 = n2164 ? wd1[10] : n1626;   // regs.v(46)
    assign n2683 = n2164 ? wd1[9] : n1627;   // regs.v(46)
    assign n2684 = n2164 ? wd1[8] : n1628;   // regs.v(46)
    assign n2685 = n2164 ? wd1[7] : n1629;   // regs.v(46)
    assign n2686 = n2164 ? wd1[6] : n1630;   // regs.v(46)
    assign n2687 = n2164 ? wd1[5] : n1631;   // regs.v(46)
    assign n2688 = n2164 ? wd1[4] : n1632;   // regs.v(46)
    assign n2689 = n2164 ? wd1[3] : n1633;   // regs.v(46)
    assign n2690 = n2164 ? wd1[2] : n1634;   // regs.v(46)
    assign n2691 = n2164 ? wd1[1] : n1635;   // regs.v(46)
    assign n2692 = n2164 ? wd1[0] : n1636;   // regs.v(46)
    assign n2693 = n2165 ? wd1[31] : n1637;   // regs.v(46)
    assign n2694 = n2165 ? wd1[30] : n1638;   // regs.v(46)
    assign n2695 = n2165 ? wd1[29] : n1639;   // regs.v(46)
    assign n2696 = n2165 ? wd1[28] : n1640;   // regs.v(46)
    assign n2697 = n2165 ? wd1[27] : n1641;   // regs.v(46)
    assign n2698 = n2165 ? wd1[26] : n1642;   // regs.v(46)
    assign n2699 = n2165 ? wd1[25] : n1643;   // regs.v(46)
    assign n2700 = n2165 ? wd1[24] : n1644;   // regs.v(46)
    assign n2701 = n2165 ? wd1[23] : n1645;   // regs.v(46)
    assign n2702 = n2165 ? wd1[22] : n1646;   // regs.v(46)
    assign n2703 = n2165 ? wd1[21] : n1647;   // regs.v(46)
    assign n2704 = n2165 ? wd1[20] : n1648;   // regs.v(46)
    assign n2705 = n2165 ? wd1[19] : n1649;   // regs.v(46)
    assign n2706 = n2165 ? wd1[18] : n1650;   // regs.v(46)
    assign n2707 = n2165 ? wd1[17] : n1651;   // regs.v(46)
    assign n2708 = n2165 ? wd1[16] : n1652;   // regs.v(46)
    assign n2709 = n2165 ? wd1[15] : n1653;   // regs.v(46)
    assign n2710 = n2165 ? wd1[14] : n1654;   // regs.v(46)
    assign n2711 = n2165 ? wd1[13] : n1655;   // regs.v(46)
    assign n2712 = n2165 ? wd1[12] : n1656;   // regs.v(46)
    assign n2713 = n2165 ? wd1[11] : n1657;   // regs.v(46)
    assign n2714 = n2165 ? wd1[10] : n1658;   // regs.v(46)
    assign n2715 = n2165 ? wd1[9] : n1659;   // regs.v(46)
    assign n2716 = n2165 ? wd1[8] : n1660;   // regs.v(46)
    assign n2717 = n2165 ? wd1[7] : n1661;   // regs.v(46)
    assign n2718 = n2165 ? wd1[6] : n1662;   // regs.v(46)
    assign n2719 = n2165 ? wd1[5] : n1663;   // regs.v(46)
    assign n2720 = n2165 ? wd1[4] : n1664;   // regs.v(46)
    assign n2721 = n2165 ? wd1[3] : n1665;   // regs.v(46)
    assign n2722 = n2165 ? wd1[2] : n1666;   // regs.v(46)
    assign n2723 = n2165 ? wd1[1] : n1667;   // regs.v(46)
    assign n2724 = n2165 ? wd1[0] : n1668;   // regs.v(46)
    assign n2725 = n2166 ? wd1[31] : n1669;   // regs.v(46)
    assign n2726 = n2166 ? wd1[30] : n1670;   // regs.v(46)
    assign n2727 = n2166 ? wd1[29] : n1671;   // regs.v(46)
    assign n2728 = n2166 ? wd1[28] : n1672;   // regs.v(46)
    assign n2729 = n2166 ? wd1[27] : n1673;   // regs.v(46)
    assign n2730 = n2166 ? wd1[26] : n1674;   // regs.v(46)
    assign n2731 = n2166 ? wd1[25] : n1675;   // regs.v(46)
    assign n2732 = n2166 ? wd1[24] : n1676;   // regs.v(46)
    assign n2733 = n2166 ? wd1[23] : n1677;   // regs.v(46)
    assign n2734 = n2166 ? wd1[22] : n1678;   // regs.v(46)
    assign n2735 = n2166 ? wd1[21] : n1679;   // regs.v(46)
    assign n2736 = n2166 ? wd1[20] : n1680;   // regs.v(46)
    assign n2737 = n2166 ? wd1[19] : n1681;   // regs.v(46)
    assign n2738 = n2166 ? wd1[18] : n1682;   // regs.v(46)
    assign n2739 = n2166 ? wd1[17] : n1683;   // regs.v(46)
    assign n2740 = n2166 ? wd1[16] : n1684;   // regs.v(46)
    assign n2741 = n2166 ? wd1[15] : n1685;   // regs.v(46)
    assign n2742 = n2166 ? wd1[14] : n1686;   // regs.v(46)
    assign n2743 = n2166 ? wd1[13] : n1687;   // regs.v(46)
    assign n2744 = n2166 ? wd1[12] : n1688;   // regs.v(46)
    assign n2745 = n2166 ? wd1[11] : n1689;   // regs.v(46)
    assign n2746 = n2166 ? wd1[10] : n1690;   // regs.v(46)
    assign n2747 = n2166 ? wd1[9] : n1691;   // regs.v(46)
    assign n2748 = n2166 ? wd1[8] : n1692;   // regs.v(46)
    assign n2749 = n2166 ? wd1[7] : n1693;   // regs.v(46)
    assign n2750 = n2166 ? wd1[6] : n1694;   // regs.v(46)
    assign n2751 = n2166 ? wd1[5] : n1695;   // regs.v(46)
    assign n2752 = n2166 ? wd1[4] : n1696;   // regs.v(46)
    assign n2753 = n2166 ? wd1[3] : n1697;   // regs.v(46)
    assign n2754 = n2166 ? wd1[2] : n1698;   // regs.v(46)
    assign n2755 = n2166 ? wd1[1] : n1699;   // regs.v(46)
    assign n2756 = n2166 ? wd1[0] : n1700;   // regs.v(46)
    assign n2757 = n2167 ? wd1[31] : n1701;   // regs.v(46)
    assign n2758 = n2167 ? wd1[30] : n1702;   // regs.v(46)
    assign n2759 = n2167 ? wd1[29] : n1703;   // regs.v(46)
    assign n2760 = n2167 ? wd1[28] : n1704;   // regs.v(46)
    assign n2761 = n2167 ? wd1[27] : n1705;   // regs.v(46)
    assign n2762 = n2167 ? wd1[26] : n1706;   // regs.v(46)
    assign n2763 = n2167 ? wd1[25] : n1707;   // regs.v(46)
    assign n2764 = n2167 ? wd1[24] : n1708;   // regs.v(46)
    assign n2765 = n2167 ? wd1[23] : n1709;   // regs.v(46)
    assign n2766 = n2167 ? wd1[22] : n1710;   // regs.v(46)
    assign n2767 = n2167 ? wd1[21] : n1711;   // regs.v(46)
    assign n2768 = n2167 ? wd1[20] : n1712;   // regs.v(46)
    assign n2769 = n2167 ? wd1[19] : n1713;   // regs.v(46)
    assign n2770 = n2167 ? wd1[18] : n1714;   // regs.v(46)
    assign n2771 = n2167 ? wd1[17] : n1715;   // regs.v(46)
    assign n2772 = n2167 ? wd1[16] : n1716;   // regs.v(46)
    assign n2773 = n2167 ? wd1[15] : n1717;   // regs.v(46)
    assign n2774 = n2167 ? wd1[14] : n1718;   // regs.v(46)
    assign n2775 = n2167 ? wd1[13] : n1719;   // regs.v(46)
    assign n2776 = n2167 ? wd1[12] : n1720;   // regs.v(46)
    assign n2777 = n2167 ? wd1[11] : n1721;   // regs.v(46)
    assign n2778 = n2167 ? wd1[10] : n1722;   // regs.v(46)
    assign n2779 = n2167 ? wd1[9] : n1723;   // regs.v(46)
    assign n2780 = n2167 ? wd1[8] : n1724;   // regs.v(46)
    assign n2781 = n2167 ? wd1[7] : n1725;   // regs.v(46)
    assign n2782 = n2167 ? wd1[6] : n1726;   // regs.v(46)
    assign n2783 = n2167 ? wd1[5] : n1727;   // regs.v(46)
    assign n2784 = n2167 ? wd1[4] : n1728;   // regs.v(46)
    assign n2785 = n2167 ? wd1[3] : n1729;   // regs.v(46)
    assign n2786 = n2167 ? wd1[2] : n1730;   // regs.v(46)
    assign n2787 = n2167 ? wd1[1] : n1731;   // regs.v(46)
    assign n2788 = n2167 ? wd1[0] : n1732;   // regs.v(46)
    assign n2789 = n2168 ? wd1[31] : n1733;   // regs.v(46)
    assign n2790 = n2168 ? wd1[30] : n1734;   // regs.v(46)
    assign n2791 = n2168 ? wd1[29] : n1735;   // regs.v(46)
    assign n2792 = n2168 ? wd1[28] : n1736;   // regs.v(46)
    assign n2793 = n2168 ? wd1[27] : n1737;   // regs.v(46)
    assign n2794 = n2168 ? wd1[26] : n1738;   // regs.v(46)
    assign n2795 = n2168 ? wd1[25] : n1739;   // regs.v(46)
    assign n2796 = n2168 ? wd1[24] : n1740;   // regs.v(46)
    assign n2797 = n2168 ? wd1[23] : n1741;   // regs.v(46)
    assign n2798 = n2168 ? wd1[22] : n1742;   // regs.v(46)
    assign n2799 = n2168 ? wd1[21] : n1743;   // regs.v(46)
    assign n2800 = n2168 ? wd1[20] : n1744;   // regs.v(46)
    assign n2801 = n2168 ? wd1[19] : n1745;   // regs.v(46)
    assign n2802 = n2168 ? wd1[18] : n1746;   // regs.v(46)
    assign n2803 = n2168 ? wd1[17] : n1747;   // regs.v(46)
    assign n2804 = n2168 ? wd1[16] : n1748;   // regs.v(46)
    assign n2805 = n2168 ? wd1[15] : n1749;   // regs.v(46)
    assign n2806 = n2168 ? wd1[14] : n1750;   // regs.v(46)
    assign n2807 = n2168 ? wd1[13] : n1751;   // regs.v(46)
    assign n2808 = n2168 ? wd1[12] : n1752;   // regs.v(46)
    assign n2809 = n2168 ? wd1[11] : n1753;   // regs.v(46)
    assign n2810 = n2168 ? wd1[10] : n1754;   // regs.v(46)
    assign n2811 = n2168 ? wd1[9] : n1755;   // regs.v(46)
    assign n2812 = n2168 ? wd1[8] : n1756;   // regs.v(46)
    assign n2813 = n2168 ? wd1[7] : n1757;   // regs.v(46)
    assign n2814 = n2168 ? wd1[6] : n1758;   // regs.v(46)
    assign n2815 = n2168 ? wd1[5] : n1759;   // regs.v(46)
    assign n2816 = n2168 ? wd1[4] : n1760;   // regs.v(46)
    assign n2817 = n2168 ? wd1[3] : n1761;   // regs.v(46)
    assign n2818 = n2168 ? wd1[2] : n1762;   // regs.v(46)
    assign n2819 = n2168 ? wd1[1] : n1763;   // regs.v(46)
    assign n2820 = n2168 ? wd1[0] : n1764;   // regs.v(46)
    assign n2821 = n2169 ? wd1[31] : n1765;   // regs.v(46)
    assign n2822 = n2169 ? wd1[30] : n1766;   // regs.v(46)
    assign n2823 = n2169 ? wd1[29] : n1767;   // regs.v(46)
    assign n2824 = n2169 ? wd1[28] : n1768;   // regs.v(46)
    assign n2825 = n2169 ? wd1[27] : n1769;   // regs.v(46)
    assign n2826 = n2169 ? wd1[26] : n1770;   // regs.v(46)
    assign n2827 = n2169 ? wd1[25] : n1771;   // regs.v(46)
    assign n2828 = n2169 ? wd1[24] : n1772;   // regs.v(46)
    assign n2829 = n2169 ? wd1[23] : n1773;   // regs.v(46)
    assign n2830 = n2169 ? wd1[22] : n1774;   // regs.v(46)
    assign n2831 = n2169 ? wd1[21] : n1775;   // regs.v(46)
    assign n2832 = n2169 ? wd1[20] : n1776;   // regs.v(46)
    assign n2833 = n2169 ? wd1[19] : n1777;   // regs.v(46)
    assign n2834 = n2169 ? wd1[18] : n1778;   // regs.v(46)
    assign n2835 = n2169 ? wd1[17] : n1779;   // regs.v(46)
    assign n2836 = n2169 ? wd1[16] : n1780;   // regs.v(46)
    assign n2837 = n2169 ? wd1[15] : n1781;   // regs.v(46)
    assign n2838 = n2169 ? wd1[14] : n1782;   // regs.v(46)
    assign n2839 = n2169 ? wd1[13] : n1783;   // regs.v(46)
    assign n2840 = n2169 ? wd1[12] : n1784;   // regs.v(46)
    assign n2841 = n2169 ? wd1[11] : n1785;   // regs.v(46)
    assign n2842 = n2169 ? wd1[10] : n1786;   // regs.v(46)
    assign n2843 = n2169 ? wd1[9] : n1787;   // regs.v(46)
    assign n2844 = n2169 ? wd1[8] : n1788;   // regs.v(46)
    assign n2845 = n2169 ? wd1[7] : n1789;   // regs.v(46)
    assign n2846 = n2169 ? wd1[6] : n1790;   // regs.v(46)
    assign n2847 = n2169 ? wd1[5] : n1791;   // regs.v(46)
    assign n2848 = n2169 ? wd1[4] : n1792;   // regs.v(46)
    assign n2849 = n2169 ? wd1[3] : n1793;   // regs.v(46)
    assign n2850 = n2169 ? wd1[2] : n1794;   // regs.v(46)
    assign n2851 = n2169 ? wd1[1] : n1795;   // regs.v(46)
    assign n2852 = n2169 ? wd1[0] : n1796;   // regs.v(46)
    assign n2853 = n2170 ? wd1[31] : n1797;   // regs.v(46)
    assign n2854 = n2170 ? wd1[30] : n1798;   // regs.v(46)
    assign n2855 = n2170 ? wd1[29] : n1799;   // regs.v(46)
    assign n2856 = n2170 ? wd1[28] : n1800;   // regs.v(46)
    assign n2857 = n2170 ? wd1[27] : n1801;   // regs.v(46)
    assign n2858 = n2170 ? wd1[26] : n1802;   // regs.v(46)
    assign n2859 = n2170 ? wd1[25] : n1803;   // regs.v(46)
    assign n2860 = n2170 ? wd1[24] : n1804;   // regs.v(46)
    assign n2861 = n2170 ? wd1[23] : n1805;   // regs.v(46)
    assign n2862 = n2170 ? wd1[22] : n1806;   // regs.v(46)
    assign n2863 = n2170 ? wd1[21] : n1807;   // regs.v(46)
    assign n2864 = n2170 ? wd1[20] : n1808;   // regs.v(46)
    assign n2865 = n2170 ? wd1[19] : n1809;   // regs.v(46)
    assign n2866 = n2170 ? wd1[18] : n1810;   // regs.v(46)
    assign n2867 = n2170 ? wd1[17] : n1811;   // regs.v(46)
    assign n2868 = n2170 ? wd1[16] : n1812;   // regs.v(46)
    assign n2869 = n2170 ? wd1[15] : n1813;   // regs.v(46)
    assign n2870 = n2170 ? wd1[14] : n1814;   // regs.v(46)
    assign n2871 = n2170 ? wd1[13] : n1815;   // regs.v(46)
    assign n2872 = n2170 ? wd1[12] : n1816;   // regs.v(46)
    assign n2873 = n2170 ? wd1[11] : n1817;   // regs.v(46)
    assign n2874 = n2170 ? wd1[10] : n1818;   // regs.v(46)
    assign n2875 = n2170 ? wd1[9] : n1819;   // regs.v(46)
    assign n2876 = n2170 ? wd1[8] : n1820;   // regs.v(46)
    assign n2877 = n2170 ? wd1[7] : n1821;   // regs.v(46)
    assign n2878 = n2170 ? wd1[6] : n1822;   // regs.v(46)
    assign n2879 = n2170 ? wd1[5] : n1823;   // regs.v(46)
    assign n2880 = n2170 ? wd1[4] : n1824;   // regs.v(46)
    assign n2881 = n2170 ? wd1[3] : n1825;   // regs.v(46)
    assign n2882 = n2170 ? wd1[2] : n1826;   // regs.v(46)
    assign n2883 = n2170 ? wd1[1] : n1827;   // regs.v(46)
    assign n2884 = n2170 ? wd1[0] : n1828;   // regs.v(46)
    assign n2885 = n2171 ? wd1[31] : n1829;   // regs.v(46)
    assign n2886 = n2171 ? wd1[30] : n1830;   // regs.v(46)
    assign n2887 = n2171 ? wd1[29] : n1831;   // regs.v(46)
    assign n2888 = n2171 ? wd1[28] : n1832;   // regs.v(46)
    assign n2889 = n2171 ? wd1[27] : n1833;   // regs.v(46)
    assign n2890 = n2171 ? wd1[26] : n1834;   // regs.v(46)
    assign n2891 = n2171 ? wd1[25] : n1835;   // regs.v(46)
    assign n2892 = n2171 ? wd1[24] : n1836;   // regs.v(46)
    assign n2893 = n2171 ? wd1[23] : n1837;   // regs.v(46)
    assign n2894 = n2171 ? wd1[22] : n1838;   // regs.v(46)
    assign n2895 = n2171 ? wd1[21] : n1839;   // regs.v(46)
    assign n2896 = n2171 ? wd1[20] : n1840;   // regs.v(46)
    assign n2897 = n2171 ? wd1[19] : n1841;   // regs.v(46)
    assign n2898 = n2171 ? wd1[18] : n1842;   // regs.v(46)
    assign n2899 = n2171 ? wd1[17] : n1843;   // regs.v(46)
    assign n2900 = n2171 ? wd1[16] : n1844;   // regs.v(46)
    assign n2901 = n2171 ? wd1[15] : n1845;   // regs.v(46)
    assign n2902 = n2171 ? wd1[14] : n1846;   // regs.v(46)
    assign n2903 = n2171 ? wd1[13] : n1847;   // regs.v(46)
    assign n2904 = n2171 ? wd1[12] : n1848;   // regs.v(46)
    assign n2905 = n2171 ? wd1[11] : n1849;   // regs.v(46)
    assign n2906 = n2171 ? wd1[10] : n1850;   // regs.v(46)
    assign n2907 = n2171 ? wd1[9] : n1851;   // regs.v(46)
    assign n2908 = n2171 ? wd1[8] : n1852;   // regs.v(46)
    assign n2909 = n2171 ? wd1[7] : n1853;   // regs.v(46)
    assign n2910 = n2171 ? wd1[6] : n1854;   // regs.v(46)
    assign n2911 = n2171 ? wd1[5] : n1855;   // regs.v(46)
    assign n2912 = n2171 ? wd1[4] : n1856;   // regs.v(46)
    assign n2913 = n2171 ? wd1[3] : n1857;   // regs.v(46)
    assign n2914 = n2171 ? wd1[2] : n1858;   // regs.v(46)
    assign n2915 = n2171 ? wd1[1] : n1859;   // regs.v(46)
    assign n2916 = n2171 ? wd1[0] : n1860;   // regs.v(46)
    assign n2917 = n2172 ? wd1[31] : n1861;   // regs.v(46)
    assign n2918 = n2172 ? wd1[30] : n1862;   // regs.v(46)
    assign n2919 = n2172 ? wd1[29] : n1863;   // regs.v(46)
    assign n2920 = n2172 ? wd1[28] : n1864;   // regs.v(46)
    assign n2921 = n2172 ? wd1[27] : n1865;   // regs.v(46)
    assign n2922 = n2172 ? wd1[26] : n1866;   // regs.v(46)
    assign n2923 = n2172 ? wd1[25] : n1867;   // regs.v(46)
    assign n2924 = n2172 ? wd1[24] : n1868;   // regs.v(46)
    assign n2925 = n2172 ? wd1[23] : n1869;   // regs.v(46)
    assign n2926 = n2172 ? wd1[22] : n1870;   // regs.v(46)
    assign n2927 = n2172 ? wd1[21] : n1871;   // regs.v(46)
    assign n2928 = n2172 ? wd1[20] : n1872;   // regs.v(46)
    assign n2929 = n2172 ? wd1[19] : n1873;   // regs.v(46)
    assign n2930 = n2172 ? wd1[18] : n1874;   // regs.v(46)
    assign n2931 = n2172 ? wd1[17] : n1875;   // regs.v(46)
    assign n2932 = n2172 ? wd1[16] : n1876;   // regs.v(46)
    assign n2933 = n2172 ? wd1[15] : n1877;   // regs.v(46)
    assign n2934 = n2172 ? wd1[14] : n1878;   // regs.v(46)
    assign n2935 = n2172 ? wd1[13] : n1879;   // regs.v(46)
    assign n2936 = n2172 ? wd1[12] : n1880;   // regs.v(46)
    assign n2937 = n2172 ? wd1[11] : n1881;   // regs.v(46)
    assign n2938 = n2172 ? wd1[10] : n1882;   // regs.v(46)
    assign n2939 = n2172 ? wd1[9] : n1883;   // regs.v(46)
    assign n2940 = n2172 ? wd1[8] : n1884;   // regs.v(46)
    assign n2941 = n2172 ? wd1[7] : n1885;   // regs.v(46)
    assign n2942 = n2172 ? wd1[6] : n1886;   // regs.v(46)
    assign n2943 = n2172 ? wd1[5] : n1887;   // regs.v(46)
    assign n2944 = n2172 ? wd1[4] : n1888;   // regs.v(46)
    assign n2945 = n2172 ? wd1[3] : n1889;   // regs.v(46)
    assign n2946 = n2172 ? wd1[2] : n1890;   // regs.v(46)
    assign n2947 = n2172 ? wd1[1] : n1891;   // regs.v(46)
    assign n2948 = n2172 ? wd1[0] : n1892;   // regs.v(46)
    assign n2949 = n2173 ? wd1[31] : n1893;   // regs.v(46)
    assign n2950 = n2173 ? wd1[30] : n1894;   // regs.v(46)
    assign n2951 = n2173 ? wd1[29] : n1895;   // regs.v(46)
    assign n2952 = n2173 ? wd1[28] : n1896;   // regs.v(46)
    assign n2953 = n2173 ? wd1[27] : n1897;   // regs.v(46)
    assign n2954 = n2173 ? wd1[26] : n1898;   // regs.v(46)
    assign n2955 = n2173 ? wd1[25] : n1899;   // regs.v(46)
    assign n2956 = n2173 ? wd1[24] : n1900;   // regs.v(46)
    assign n2957 = n2173 ? wd1[23] : n1901;   // regs.v(46)
    assign n2958 = n2173 ? wd1[22] : n1902;   // regs.v(46)
    assign n2959 = n2173 ? wd1[21] : n1903;   // regs.v(46)
    assign n2960 = n2173 ? wd1[20] : n1904;   // regs.v(46)
    assign n2961 = n2173 ? wd1[19] : n1905;   // regs.v(46)
    assign n2962 = n2173 ? wd1[18] : n1906;   // regs.v(46)
    assign n2963 = n2173 ? wd1[17] : n1907;   // regs.v(46)
    assign n2964 = n2173 ? wd1[16] : n1908;   // regs.v(46)
    assign n2965 = n2173 ? wd1[15] : n1909;   // regs.v(46)
    assign n2966 = n2173 ? wd1[14] : n1910;   // regs.v(46)
    assign n2967 = n2173 ? wd1[13] : n1911;   // regs.v(46)
    assign n2968 = n2173 ? wd1[12] : n1912;   // regs.v(46)
    assign n2969 = n2173 ? wd1[11] : n1913;   // regs.v(46)
    assign n2970 = n2173 ? wd1[10] : n1914;   // regs.v(46)
    assign n2971 = n2173 ? wd1[9] : n1915;   // regs.v(46)
    assign n2972 = n2173 ? wd1[8] : n1916;   // regs.v(46)
    assign n2973 = n2173 ? wd1[7] : n1917;   // regs.v(46)
    assign n2974 = n2173 ? wd1[6] : n1918;   // regs.v(46)
    assign n2975 = n2173 ? wd1[5] : n1919;   // regs.v(46)
    assign n2976 = n2173 ? wd1[4] : n1920;   // regs.v(46)
    assign n2977 = n2173 ? wd1[3] : n1921;   // regs.v(46)
    assign n2978 = n2173 ? wd1[2] : n1922;   // regs.v(46)
    assign n2979 = n2173 ? wd1[1] : n1923;   // regs.v(46)
    assign n2980 = n2173 ? wd1[0] : n1924;   // regs.v(46)
    assign n2981 = n2174 ? wd1[31] : n1925;   // regs.v(46)
    assign n2982 = n2174 ? wd1[30] : n1926;   // regs.v(46)
    assign n2983 = n2174 ? wd1[29] : n1927;   // regs.v(46)
    assign n2984 = n2174 ? wd1[28] : n1928;   // regs.v(46)
    assign n2985 = n2174 ? wd1[27] : n1929;   // regs.v(46)
    assign n2986 = n2174 ? wd1[26] : n1930;   // regs.v(46)
    assign n2987 = n2174 ? wd1[25] : n1931;   // regs.v(46)
    assign n2988 = n2174 ? wd1[24] : n1932;   // regs.v(46)
    assign n2989 = n2174 ? wd1[23] : n1933;   // regs.v(46)
    assign n2990 = n2174 ? wd1[22] : n1934;   // regs.v(46)
    assign n2991 = n2174 ? wd1[21] : n1935;   // regs.v(46)
    assign n2992 = n2174 ? wd1[20] : n1936;   // regs.v(46)
    assign n2993 = n2174 ? wd1[19] : n1937;   // regs.v(46)
    assign n2994 = n2174 ? wd1[18] : n1938;   // regs.v(46)
    assign n2995 = n2174 ? wd1[17] : n1939;   // regs.v(46)
    assign n2996 = n2174 ? wd1[16] : n1940;   // regs.v(46)
    assign n2997 = n2174 ? wd1[15] : n1941;   // regs.v(46)
    assign n2998 = n2174 ? wd1[14] : n1942;   // regs.v(46)
    assign n2999 = n2174 ? wd1[13] : n1943;   // regs.v(46)
    assign n3000 = n2174 ? wd1[12] : n1944;   // regs.v(46)
    assign n3001 = n2174 ? wd1[11] : n1945;   // regs.v(46)
    assign n3002 = n2174 ? wd1[10] : n1946;   // regs.v(46)
    assign n3003 = n2174 ? wd1[9] : n1947;   // regs.v(46)
    assign n3004 = n2174 ? wd1[8] : n1948;   // regs.v(46)
    assign n3005 = n2174 ? wd1[7] : n1949;   // regs.v(46)
    assign n3006 = n2174 ? wd1[6] : n1950;   // regs.v(46)
    assign n3007 = n2174 ? wd1[5] : n1951;   // regs.v(46)
    assign n3008 = n2174 ? wd1[4] : n1952;   // regs.v(46)
    assign n3009 = n2174 ? wd1[3] : n1953;   // regs.v(46)
    assign n3010 = n2174 ? wd1[2] : n1954;   // regs.v(46)
    assign n3011 = n2174 ? wd1[1] : n1955;   // regs.v(46)
    assign n3012 = n2174 ? wd1[0] : n1956;   // regs.v(46)
    assign n3013 = n2175 ? wd1[31] : n1957;   // regs.v(46)
    assign n3014 = n2175 ? wd1[30] : n1958;   // regs.v(46)
    assign n3015 = n2175 ? wd1[29] : n1959;   // regs.v(46)
    assign n3016 = n2175 ? wd1[28] : n1960;   // regs.v(46)
    assign n3017 = n2175 ? wd1[27] : n1961;   // regs.v(46)
    assign n3018 = n2175 ? wd1[26] : n1962;   // regs.v(46)
    assign n3019 = n2175 ? wd1[25] : n1963;   // regs.v(46)
    assign n3020 = n2175 ? wd1[24] : n1964;   // regs.v(46)
    assign n3021 = n2175 ? wd1[23] : n1965;   // regs.v(46)
    assign n3022 = n2175 ? wd1[22] : n1966;   // regs.v(46)
    assign n3023 = n2175 ? wd1[21] : n1967;   // regs.v(46)
    assign n3024 = n2175 ? wd1[20] : n1968;   // regs.v(46)
    assign n3025 = n2175 ? wd1[19] : n1969;   // regs.v(46)
    assign n3026 = n2175 ? wd1[18] : n1970;   // regs.v(46)
    assign n3027 = n2175 ? wd1[17] : n1971;   // regs.v(46)
    assign n3028 = n2175 ? wd1[16] : n1972;   // regs.v(46)
    assign n3029 = n2175 ? wd1[15] : n1973;   // regs.v(46)
    assign n3030 = n2175 ? wd1[14] : n1974;   // regs.v(46)
    assign n3031 = n2175 ? wd1[13] : n1975;   // regs.v(46)
    assign n3032 = n2175 ? wd1[12] : n1976;   // regs.v(46)
    assign n3033 = n2175 ? wd1[11] : n1977;   // regs.v(46)
    assign n3034 = n2175 ? wd1[10] : n1978;   // regs.v(46)
    assign n3035 = n2175 ? wd1[9] : n1979;   // regs.v(46)
    assign n3036 = n2175 ? wd1[8] : n1980;   // regs.v(46)
    assign n3037 = n2175 ? wd1[7] : n1981;   // regs.v(46)
    assign n3038 = n2175 ? wd1[6] : n1982;   // regs.v(46)
    assign n3039 = n2175 ? wd1[5] : n1983;   // regs.v(46)
    assign n3040 = n2175 ? wd1[4] : n1984;   // regs.v(46)
    assign n3041 = n2175 ? wd1[3] : n1985;   // regs.v(46)
    assign n3042 = n2175 ? wd1[2] : n1986;   // regs.v(46)
    assign n3043 = n2175 ? wd1[1] : n1987;   // regs.v(46)
    assign n3044 = n2175 ? wd1[0] : n1988;   // regs.v(46)
    assign n3045 = n2176 ? wd1[31] : n1989;   // regs.v(46)
    assign n3046 = n2176 ? wd1[30] : n1990;   // regs.v(46)
    assign n3047 = n2176 ? wd1[29] : n1991;   // regs.v(46)
    assign n3048 = n2176 ? wd1[28] : n1992;   // regs.v(46)
    assign n3049 = n2176 ? wd1[27] : n1993;   // regs.v(46)
    assign n3050 = n2176 ? wd1[26] : n1994;   // regs.v(46)
    assign n3051 = n2176 ? wd1[25] : n1995;   // regs.v(46)
    assign n3052 = n2176 ? wd1[24] : n1996;   // regs.v(46)
    assign n3053 = n2176 ? wd1[23] : n1997;   // regs.v(46)
    assign n3054 = n2176 ? wd1[22] : n1998;   // regs.v(46)
    assign n3055 = n2176 ? wd1[21] : n1999;   // regs.v(46)
    assign n3056 = n2176 ? wd1[20] : n2000;   // regs.v(46)
    assign n3057 = n2176 ? wd1[19] : n2001;   // regs.v(46)
    assign n3058 = n2176 ? wd1[18] : n2002;   // regs.v(46)
    assign n3059 = n2176 ? wd1[17] : n2003;   // regs.v(46)
    assign n3060 = n2176 ? wd1[16] : n2004;   // regs.v(46)
    assign n3061 = n2176 ? wd1[15] : n2005;   // regs.v(46)
    assign n3062 = n2176 ? wd1[14] : n2006;   // regs.v(46)
    assign n3063 = n2176 ? wd1[13] : n2007;   // regs.v(46)
    assign n3064 = n2176 ? wd1[12] : n2008;   // regs.v(46)
    assign n3065 = n2176 ? wd1[11] : n2009;   // regs.v(46)
    assign n3066 = n2176 ? wd1[10] : n2010;   // regs.v(46)
    assign n3067 = n2176 ? wd1[9] : n2011;   // regs.v(46)
    assign n3068 = n2176 ? wd1[8] : n2012;   // regs.v(46)
    assign n3069 = n2176 ? wd1[7] : n2013;   // regs.v(46)
    assign n3070 = n2176 ? wd1[6] : n2014;   // regs.v(46)
    assign n3071 = n2176 ? wd1[5] : n2015;   // regs.v(46)
    assign n3072 = n2176 ? wd1[4] : n2016;   // regs.v(46)
    assign n3073 = n2176 ? wd1[3] : n2017;   // regs.v(46)
    assign n3074 = n2176 ? wd1[2] : n2018;   // regs.v(46)
    assign n3075 = n2176 ? wd1[1] : n2019;   // regs.v(46)
    assign n3076 = n2176 ? wd1[0] : n2020;   // regs.v(46)
    assign n3077 = n2177 ? wd1[31] : n2021;   // regs.v(46)
    assign n3078 = n2177 ? wd1[30] : n2022;   // regs.v(46)
    assign n3079 = n2177 ? wd1[29] : n2023;   // regs.v(46)
    assign n3080 = n2177 ? wd1[28] : n2024;   // regs.v(46)
    assign n3081 = n2177 ? wd1[27] : n2025;   // regs.v(46)
    assign n3082 = n2177 ? wd1[26] : n2026;   // regs.v(46)
    assign n3083 = n2177 ? wd1[25] : n2027;   // regs.v(46)
    assign n3084 = n2177 ? wd1[24] : n2028;   // regs.v(46)
    assign n3085 = n2177 ? wd1[23] : n2029;   // regs.v(46)
    assign n3086 = n2177 ? wd1[22] : n2030;   // regs.v(46)
    assign n3087 = n2177 ? wd1[21] : n2031;   // regs.v(46)
    assign n3088 = n2177 ? wd1[20] : n2032;   // regs.v(46)
    assign n3089 = n2177 ? wd1[19] : n2033;   // regs.v(46)
    assign n3090 = n2177 ? wd1[18] : n2034;   // regs.v(46)
    assign n3091 = n2177 ? wd1[17] : n2035;   // regs.v(46)
    assign n3092 = n2177 ? wd1[16] : n2036;   // regs.v(46)
    assign n3093 = n2177 ? wd1[15] : n2037;   // regs.v(46)
    assign n3094 = n2177 ? wd1[14] : n2038;   // regs.v(46)
    assign n3095 = n2177 ? wd1[13] : n2039;   // regs.v(46)
    assign n3096 = n2177 ? wd1[12] : n2040;   // regs.v(46)
    assign n3097 = n2177 ? wd1[11] : n2041;   // regs.v(46)
    assign n3098 = n2177 ? wd1[10] : n2042;   // regs.v(46)
    assign n3099 = n2177 ? wd1[9] : n2043;   // regs.v(46)
    assign n3100 = n2177 ? wd1[8] : n2044;   // regs.v(46)
    assign n3101 = n2177 ? wd1[7] : n2045;   // regs.v(46)
    assign n3102 = n2177 ? wd1[6] : n2046;   // regs.v(46)
    assign n3103 = n2177 ? wd1[5] : n2047;   // regs.v(46)
    assign n3104 = n2177 ? wd1[4] : n2048;   // regs.v(46)
    assign n3105 = n2177 ? wd1[3] : n2049;   // regs.v(46)
    assign n3106 = n2177 ? wd1[2] : n2050;   // regs.v(46)
    assign n3107 = n2177 ? wd1[1] : n2051;   // regs.v(46)
    assign n3108 = n2177 ? wd1[0] : n2052;   // regs.v(46)
    assign n3109 = n2178 ? wd1[31] : n2053;   // regs.v(46)
    assign n3110 = n2178 ? wd1[30] : n2054;   // regs.v(46)
    assign n3111 = n2178 ? wd1[29] : n2055;   // regs.v(46)
    assign n3112 = n2178 ? wd1[28] : n2056;   // regs.v(46)
    assign n3113 = n2178 ? wd1[27] : n2057;   // regs.v(46)
    assign n3114 = n2178 ? wd1[26] : n2058;   // regs.v(46)
    assign n3115 = n2178 ? wd1[25] : n2059;   // regs.v(46)
    assign n3116 = n2178 ? wd1[24] : n2060;   // regs.v(46)
    assign n3117 = n2178 ? wd1[23] : n2061;   // regs.v(46)
    assign n3118 = n2178 ? wd1[22] : n2062;   // regs.v(46)
    assign n3119 = n2178 ? wd1[21] : n2063;   // regs.v(46)
    assign n3120 = n2178 ? wd1[20] : n2064;   // regs.v(46)
    assign n3121 = n2178 ? wd1[19] : n2065;   // regs.v(46)
    assign n3122 = n2178 ? wd1[18] : n2066;   // regs.v(46)
    assign n3123 = n2178 ? wd1[17] : n2067;   // regs.v(46)
    assign n3124 = n2178 ? wd1[16] : n2068;   // regs.v(46)
    assign n3125 = n2178 ? wd1[15] : n2069;   // regs.v(46)
    assign n3126 = n2178 ? wd1[14] : n2070;   // regs.v(46)
    assign n3127 = n2178 ? wd1[13] : n2071;   // regs.v(46)
    assign n3128 = n2178 ? wd1[12] : n2072;   // regs.v(46)
    assign n3129 = n2178 ? wd1[11] : n2073;   // regs.v(46)
    assign n3130 = n2178 ? wd1[10] : n2074;   // regs.v(46)
    assign n3131 = n2178 ? wd1[9] : n2075;   // regs.v(46)
    assign n3132 = n2178 ? wd1[8] : n2076;   // regs.v(46)
    assign n3133 = n2178 ? wd1[7] : n2077;   // regs.v(46)
    assign n3134 = n2178 ? wd1[6] : n2078;   // regs.v(46)
    assign n3135 = n2178 ? wd1[5] : n2079;   // regs.v(46)
    assign n3136 = n2178 ? wd1[4] : n2080;   // regs.v(46)
    assign n3137 = n2178 ? wd1[3] : n2081;   // regs.v(46)
    assign n3138 = n2178 ? wd1[2] : n2082;   // regs.v(46)
    assign n3139 = n2178 ? wd1[1] : n2083;   // regs.v(46)
    assign n3140 = n2178 ? wd1[0] : n2084;   // regs.v(46)
    assign n3141 = n2179 ? wd1[31] : n2085;   // regs.v(46)
    assign n3142 = n2179 ? wd1[30] : n2086;   // regs.v(46)
    assign n3143 = n2179 ? wd1[29] : n2087;   // regs.v(46)
    assign n3144 = n2179 ? wd1[28] : n2088;   // regs.v(46)
    assign n3145 = n2179 ? wd1[27] : n2089;   // regs.v(46)
    assign n3146 = n2179 ? wd1[26] : n2090;   // regs.v(46)
    assign n3147 = n2179 ? wd1[25] : n2091;   // regs.v(46)
    assign n3148 = n2179 ? wd1[24] : n2092;   // regs.v(46)
    assign n3149 = n2179 ? wd1[23] : n2093;   // regs.v(46)
    assign n3150 = n2179 ? wd1[22] : n2094;   // regs.v(46)
    assign n3151 = n2179 ? wd1[21] : n2095;   // regs.v(46)
    assign n3152 = n2179 ? wd1[20] : n2096;   // regs.v(46)
    assign n3153 = n2179 ? wd1[19] : n2097;   // regs.v(46)
    assign n3154 = n2179 ? wd1[18] : n2098;   // regs.v(46)
    assign n3155 = n2179 ? wd1[17] : n2099;   // regs.v(46)
    assign n3156 = n2179 ? wd1[16] : n2100;   // regs.v(46)
    assign n3157 = n2179 ? wd1[15] : n2101;   // regs.v(46)
    assign n3158 = n2179 ? wd1[14] : n2102;   // regs.v(46)
    assign n3159 = n2179 ? wd1[13] : n2103;   // regs.v(46)
    assign n3160 = n2179 ? wd1[12] : n2104;   // regs.v(46)
    assign n3161 = n2179 ? wd1[11] : n2105;   // regs.v(46)
    assign n3162 = n2179 ? wd1[10] : n2106;   // regs.v(46)
    assign n3163 = n2179 ? wd1[9] : n2107;   // regs.v(46)
    assign n3164 = n2179 ? wd1[8] : n2108;   // regs.v(46)
    assign n3165 = n2179 ? wd1[7] : n2109;   // regs.v(46)
    assign n3166 = n2179 ? wd1[6] : n2110;   // regs.v(46)
    assign n3167 = n2179 ? wd1[5] : n2111;   // regs.v(46)
    assign n3168 = n2179 ? wd1[4] : n2112;   // regs.v(46)
    assign n3169 = n2179 ? wd1[3] : n2113;   // regs.v(46)
    assign n3170 = n2179 ? wd1[2] : n2114;   // regs.v(46)
    assign n3171 = n2179 ? wd1[1] : n2115;   // regs.v(46)
    assign n3172 = n2179 ? wd1[0] : n2116;   // regs.v(46)
    assign n3173 = n2180 ? wd1[31] : n2117;   // regs.v(46)
    assign n3174 = n2180 ? wd1[30] : n2118;   // regs.v(46)
    assign n3175 = n2180 ? wd1[29] : n2119;   // regs.v(46)
    assign n3176 = n2180 ? wd1[28] : n2120;   // regs.v(46)
    assign n3177 = n2180 ? wd1[27] : n2121;   // regs.v(46)
    assign n3178 = n2180 ? wd1[26] : n2122;   // regs.v(46)
    assign n3179 = n2180 ? wd1[25] : n2123;   // regs.v(46)
    assign n3180 = n2180 ? wd1[24] : n2124;   // regs.v(46)
    assign n3181 = n2180 ? wd1[23] : n2125;   // regs.v(46)
    assign n3182 = n2180 ? wd1[22] : n2126;   // regs.v(46)
    assign n3183 = n2180 ? wd1[21] : n2127;   // regs.v(46)
    assign n3184 = n2180 ? wd1[20] : n2128;   // regs.v(46)
    assign n3185 = n2180 ? wd1[19] : n2129;   // regs.v(46)
    assign n3186 = n2180 ? wd1[18] : n2130;   // regs.v(46)
    assign n3187 = n2180 ? wd1[17] : n2131;   // regs.v(46)
    assign n3188 = n2180 ? wd1[16] : n2132;   // regs.v(46)
    assign n3189 = n2180 ? wd1[15] : n2133;   // regs.v(46)
    assign n3190 = n2180 ? wd1[14] : n2134;   // regs.v(46)
    assign n3191 = n2180 ? wd1[13] : n2135;   // regs.v(46)
    assign n3192 = n2180 ? wd1[12] : n2136;   // regs.v(46)
    assign n3193 = n2180 ? wd1[11] : n2137;   // regs.v(46)
    assign n3194 = n2180 ? wd1[10] : n2138;   // regs.v(46)
    assign n3195 = n2180 ? wd1[9] : n2139;   // regs.v(46)
    assign n3196 = n2180 ? wd1[8] : n2140;   // regs.v(46)
    assign n3197 = n2180 ? wd1[7] : n2141;   // regs.v(46)
    assign n3198 = n2180 ? wd1[6] : n2142;   // regs.v(46)
    assign n3199 = n2180 ? wd1[5] : n2143;   // regs.v(46)
    assign n3200 = n2180 ? wd1[4] : n2144;   // regs.v(46)
    assign n3201 = n2180 ? wd1[3] : n2145;   // regs.v(46)
    assign n3202 = n2180 ? wd1[2] : n2146;   // regs.v(46)
    assign n3203 = n2180 ? wd1[1] : n2147;   // regs.v(46)
    assign n3204 = n2180 ? wd1[0] : n2148;   // regs.v(46)
    assign n3205 = write[1] ? n2181 : n1125;   // regs.v(46)
    assign n3206 = write[1] ? n2182 : n1126;   // regs.v(46)
    assign n3207 = write[1] ? n2183 : n1127;   // regs.v(46)
    assign n3208 = write[1] ? n2184 : n1128;   // regs.v(46)
    assign n3209 = write[1] ? n2185 : n1129;   // regs.v(46)
    assign n3210 = write[1] ? n2186 : n1130;   // regs.v(46)
    assign n3211 = write[1] ? n2187 : n1131;   // regs.v(46)
    assign n3212 = write[1] ? n2188 : n1132;   // regs.v(46)
    assign n3213 = write[1] ? n2189 : n1133;   // regs.v(46)
    assign n3214 = write[1] ? n2190 : n1134;   // regs.v(46)
    assign n3215 = write[1] ? n2191 : n1135;   // regs.v(46)
    assign n3216 = write[1] ? n2192 : n1136;   // regs.v(46)
    assign n3217 = write[1] ? n2193 : n1137;   // regs.v(46)
    assign n3218 = write[1] ? n2194 : n1138;   // regs.v(46)
    assign n3219 = write[1] ? n2195 : n1139;   // regs.v(46)
    assign n3220 = write[1] ? n2196 : n1140;   // regs.v(46)
    assign n3221 = write[1] ? n2197 : n1141;   // regs.v(46)
    assign n3222 = write[1] ? n2198 : n1142;   // regs.v(46)
    assign n3223 = write[1] ? n2199 : n1143;   // regs.v(46)
    assign n3224 = write[1] ? n2200 : n1144;   // regs.v(46)
    assign n3225 = write[1] ? n2201 : n1145;   // regs.v(46)
    assign n3226 = write[1] ? n2202 : n1146;   // regs.v(46)
    assign n3227 = write[1] ? n2203 : n1147;   // regs.v(46)
    assign n3228 = write[1] ? n2204 : n1148;   // regs.v(46)
    assign n3229 = write[1] ? n2205 : n1149;   // regs.v(46)
    assign n3230 = write[1] ? n2206 : n1150;   // regs.v(46)
    assign n3231 = write[1] ? n2207 : n1151;   // regs.v(46)
    assign n3232 = write[1] ? n2208 : n1152;   // regs.v(46)
    assign n3233 = write[1] ? n2209 : n1153;   // regs.v(46)
    assign n3234 = write[1] ? n2210 : n1154;   // regs.v(46)
    assign n3235 = write[1] ? n2211 : n1155;   // regs.v(46)
    assign n3236 = write[1] ? n2212 : n1156;   // regs.v(46)
    assign n3237 = write[1] ? n2213 : n1157;   // regs.v(46)
    assign n3238 = write[1] ? n2214 : n1158;   // regs.v(46)
    assign n3239 = write[1] ? n2215 : n1159;   // regs.v(46)
    assign n3240 = write[1] ? n2216 : n1160;   // regs.v(46)
    assign n3241 = write[1] ? n2217 : n1161;   // regs.v(46)
    assign n3242 = write[1] ? n2218 : n1162;   // regs.v(46)
    assign n3243 = write[1] ? n2219 : n1163;   // regs.v(46)
    assign n3244 = write[1] ? n2220 : n1164;   // regs.v(46)
    assign n3245 = write[1] ? n2221 : n1165;   // regs.v(46)
    assign n3246 = write[1] ? n2222 : n1166;   // regs.v(46)
    assign n3247 = write[1] ? n2223 : n1167;   // regs.v(46)
    assign n3248 = write[1] ? n2224 : n1168;   // regs.v(46)
    assign n3249 = write[1] ? n2225 : n1169;   // regs.v(46)
    assign n3250 = write[1] ? n2226 : n1170;   // regs.v(46)
    assign n3251 = write[1] ? n2227 : n1171;   // regs.v(46)
    assign n3252 = write[1] ? n2228 : n1172;   // regs.v(46)
    assign n3253 = write[1] ? n2229 : n1173;   // regs.v(46)
    assign n3254 = write[1] ? n2230 : n1174;   // regs.v(46)
    assign n3255 = write[1] ? n2231 : n1175;   // regs.v(46)
    assign n3256 = write[1] ? n2232 : n1176;   // regs.v(46)
    assign n3257 = write[1] ? n2233 : n1177;   // regs.v(46)
    assign n3258 = write[1] ? n2234 : n1178;   // regs.v(46)
    assign n3259 = write[1] ? n2235 : n1179;   // regs.v(46)
    assign n3260 = write[1] ? n2236 : n1180;   // regs.v(46)
    assign n3261 = write[1] ? n2237 : n1181;   // regs.v(46)
    assign n3262 = write[1] ? n2238 : n1182;   // regs.v(46)
    assign n3263 = write[1] ? n2239 : n1183;   // regs.v(46)
    assign n3264 = write[1] ? n2240 : n1184;   // regs.v(46)
    assign n3265 = write[1] ? n2241 : n1185;   // regs.v(46)
    assign n3266 = write[1] ? n2242 : n1186;   // regs.v(46)
    assign n3267 = write[1] ? n2243 : n1187;   // regs.v(46)
    assign n3268 = write[1] ? n2244 : n1188;   // regs.v(46)
    assign n3269 = write[1] ? n2245 : n1189;   // regs.v(46)
    assign n3270 = write[1] ? n2246 : n1190;   // regs.v(46)
    assign n3271 = write[1] ? n2247 : n1191;   // regs.v(46)
    assign n3272 = write[1] ? n2248 : n1192;   // regs.v(46)
    assign n3273 = write[1] ? n2249 : n1193;   // regs.v(46)
    assign n3274 = write[1] ? n2250 : n1194;   // regs.v(46)
    assign n3275 = write[1] ? n2251 : n1195;   // regs.v(46)
    assign n3276 = write[1] ? n2252 : n1196;   // regs.v(46)
    assign n3277 = write[1] ? n2253 : n1197;   // regs.v(46)
    assign n3278 = write[1] ? n2254 : n1198;   // regs.v(46)
    assign n3279 = write[1] ? n2255 : n1199;   // regs.v(46)
    assign n3280 = write[1] ? n2256 : n1200;   // regs.v(46)
    assign n3281 = write[1] ? n2257 : n1201;   // regs.v(46)
    assign n3282 = write[1] ? n2258 : n1202;   // regs.v(46)
    assign n3283 = write[1] ? n2259 : n1203;   // regs.v(46)
    assign n3284 = write[1] ? n2260 : n1204;   // regs.v(46)
    assign n3285 = write[1] ? n2261 : n1205;   // regs.v(46)
    assign n3286 = write[1] ? n2262 : n1206;   // regs.v(46)
    assign n3287 = write[1] ? n2263 : n1207;   // regs.v(46)
    assign n3288 = write[1] ? n2264 : n1208;   // regs.v(46)
    assign n3289 = write[1] ? n2265 : n1209;   // regs.v(46)
    assign n3290 = write[1] ? n2266 : n1210;   // regs.v(46)
    assign n3291 = write[1] ? n2267 : n1211;   // regs.v(46)
    assign n3292 = write[1] ? n2268 : n1212;   // regs.v(46)
    assign n3293 = write[1] ? n2269 : n1213;   // regs.v(46)
    assign n3294 = write[1] ? n2270 : n1214;   // regs.v(46)
    assign n3295 = write[1] ? n2271 : n1215;   // regs.v(46)
    assign n3296 = write[1] ? n2272 : n1216;   // regs.v(46)
    assign n3297 = write[1] ? n2273 : n1217;   // regs.v(46)
    assign n3298 = write[1] ? n2274 : n1218;   // regs.v(46)
    assign n3299 = write[1] ? n2275 : n1219;   // regs.v(46)
    assign n3300 = write[1] ? n2276 : n1220;   // regs.v(46)
    assign n3301 = write[1] ? n2277 : n1221;   // regs.v(46)
    assign n3302 = write[1] ? n2278 : n1222;   // regs.v(46)
    assign n3303 = write[1] ? n2279 : n1223;   // regs.v(46)
    assign n3304 = write[1] ? n2280 : n1224;   // regs.v(46)
    assign n3305 = write[1] ? n2281 : n1225;   // regs.v(46)
    assign n3306 = write[1] ? n2282 : n1226;   // regs.v(46)
    assign n3307 = write[1] ? n2283 : n1227;   // regs.v(46)
    assign n3308 = write[1] ? n2284 : n1228;   // regs.v(46)
    assign n3309 = write[1] ? n2285 : n1229;   // regs.v(46)
    assign n3310 = write[1] ? n2286 : n1230;   // regs.v(46)
    assign n3311 = write[1] ? n2287 : n1231;   // regs.v(46)
    assign n3312 = write[1] ? n2288 : n1232;   // regs.v(46)
    assign n3313 = write[1] ? n2289 : n1233;   // regs.v(46)
    assign n3314 = write[1] ? n2290 : n1234;   // regs.v(46)
    assign n3315 = write[1] ? n2291 : n1235;   // regs.v(46)
    assign n3316 = write[1] ? n2292 : n1236;   // regs.v(46)
    assign n3317 = write[1] ? n2293 : n1237;   // regs.v(46)
    assign n3318 = write[1] ? n2294 : n1238;   // regs.v(46)
    assign n3319 = write[1] ? n2295 : n1239;   // regs.v(46)
    assign n3320 = write[1] ? n2296 : n1240;   // regs.v(46)
    assign n3321 = write[1] ? n2297 : n1241;   // regs.v(46)
    assign n3322 = write[1] ? n2298 : n1242;   // regs.v(46)
    assign n3323 = write[1] ? n2299 : n1243;   // regs.v(46)
    assign n3324 = write[1] ? n2300 : n1244;   // regs.v(46)
    assign n3325 = write[1] ? n2301 : n1245;   // regs.v(46)
    assign n3326 = write[1] ? n2302 : n1246;   // regs.v(46)
    assign n3327 = write[1] ? n2303 : n1247;   // regs.v(46)
    assign n3328 = write[1] ? n2304 : n1248;   // regs.v(46)
    assign n3329 = write[1] ? n2305 : n1249;   // regs.v(46)
    assign n3330 = write[1] ? n2306 : n1250;   // regs.v(46)
    assign n3331 = write[1] ? n2307 : n1251;   // regs.v(46)
    assign n3332 = write[1] ? n2308 : n1252;   // regs.v(46)
    assign n3333 = write[1] ? n2309 : n1253;   // regs.v(46)
    assign n3334 = write[1] ? n2310 : n1254;   // regs.v(46)
    assign n3335 = write[1] ? n2311 : n1255;   // regs.v(46)
    assign n3336 = write[1] ? n2312 : n1256;   // regs.v(46)
    assign n3337 = write[1] ? n2313 : n1257;   // regs.v(46)
    assign n3338 = write[1] ? n2314 : n1258;   // regs.v(46)
    assign n3339 = write[1] ? n2315 : n1259;   // regs.v(46)
    assign n3340 = write[1] ? n2316 : n1260;   // regs.v(46)
    assign n3341 = write[1] ? n2317 : n1261;   // regs.v(46)
    assign n3342 = write[1] ? n2318 : n1262;   // regs.v(46)
    assign n3343 = write[1] ? n2319 : n1263;   // regs.v(46)
    assign n3344 = write[1] ? n2320 : n1264;   // regs.v(46)
    assign n3345 = write[1] ? n2321 : n1265;   // regs.v(46)
    assign n3346 = write[1] ? n2322 : n1266;   // regs.v(46)
    assign n3347 = write[1] ? n2323 : n1267;   // regs.v(46)
    assign n3348 = write[1] ? n2324 : n1268;   // regs.v(46)
    assign n3349 = write[1] ? n2325 : n1269;   // regs.v(46)
    assign n3350 = write[1] ? n2326 : n1270;   // regs.v(46)
    assign n3351 = write[1] ? n2327 : n1271;   // regs.v(46)
    assign n3352 = write[1] ? n2328 : n1272;   // regs.v(46)
    assign n3353 = write[1] ? n2329 : n1273;   // regs.v(46)
    assign n3354 = write[1] ? n2330 : n1274;   // regs.v(46)
    assign n3355 = write[1] ? n2331 : n1275;   // regs.v(46)
    assign n3356 = write[1] ? n2332 : n1276;   // regs.v(46)
    assign n3357 = write[1] ? n2333 : n1277;   // regs.v(46)
    assign n3358 = write[1] ? n2334 : n1278;   // regs.v(46)
    assign n3359 = write[1] ? n2335 : n1279;   // regs.v(46)
    assign n3360 = write[1] ? n2336 : n1280;   // regs.v(46)
    assign n3361 = write[1] ? n2337 : n1281;   // regs.v(46)
    assign n3362 = write[1] ? n2338 : n1282;   // regs.v(46)
    assign n3363 = write[1] ? n2339 : n1283;   // regs.v(46)
    assign n3364 = write[1] ? n2340 : n1284;   // regs.v(46)
    assign n3365 = write[1] ? n2341 : n1285;   // regs.v(46)
    assign n3366 = write[1] ? n2342 : n1286;   // regs.v(46)
    assign n3367 = write[1] ? n2343 : n1287;   // regs.v(46)
    assign n3368 = write[1] ? n2344 : n1288;   // regs.v(46)
    assign n3369 = write[1] ? n2345 : n1289;   // regs.v(46)
    assign n3370 = write[1] ? n2346 : n1290;   // regs.v(46)
    assign n3371 = write[1] ? n2347 : n1291;   // regs.v(46)
    assign n3372 = write[1] ? n2348 : n1292;   // regs.v(46)
    assign n3373 = write[1] ? n2349 : n1293;   // regs.v(46)
    assign n3374 = write[1] ? n2350 : n1294;   // regs.v(46)
    assign n3375 = write[1] ? n2351 : n1295;   // regs.v(46)
    assign n3376 = write[1] ? n2352 : n1296;   // regs.v(46)
    assign n3377 = write[1] ? n2353 : n1297;   // regs.v(46)
    assign n3378 = write[1] ? n2354 : n1298;   // regs.v(46)
    assign n3379 = write[1] ? n2355 : n1299;   // regs.v(46)
    assign n3380 = write[1] ? n2356 : n1300;   // regs.v(46)
    assign n3381 = write[1] ? n2357 : n1301;   // regs.v(46)
    assign n3382 = write[1] ? n2358 : n1302;   // regs.v(46)
    assign n3383 = write[1] ? n2359 : n1303;   // regs.v(46)
    assign n3384 = write[1] ? n2360 : n1304;   // regs.v(46)
    assign n3385 = write[1] ? n2361 : n1305;   // regs.v(46)
    assign n3386 = write[1] ? n2362 : n1306;   // regs.v(46)
    assign n3387 = write[1] ? n2363 : n1307;   // regs.v(46)
    assign n3388 = write[1] ? n2364 : n1308;   // regs.v(46)
    assign n3389 = write[1] ? n2365 : n1309;   // regs.v(46)
    assign n3390 = write[1] ? n2366 : n1310;   // regs.v(46)
    assign n3391 = write[1] ? n2367 : n1311;   // regs.v(46)
    assign n3392 = write[1] ? n2368 : n1312;   // regs.v(46)
    assign n3393 = write[1] ? n2369 : n1313;   // regs.v(46)
    assign n3394 = write[1] ? n2370 : n1314;   // regs.v(46)
    assign n3395 = write[1] ? n2371 : n1315;   // regs.v(46)
    assign n3396 = write[1] ? n2372 : n1316;   // regs.v(46)
    assign n3397 = write[1] ? n2373 : n1317;   // regs.v(46)
    assign n3398 = write[1] ? n2374 : n1318;   // regs.v(46)
    assign n3399 = write[1] ? n2375 : n1319;   // regs.v(46)
    assign n3400 = write[1] ? n2376 : n1320;   // regs.v(46)
    assign n3401 = write[1] ? n2377 : n1321;   // regs.v(46)
    assign n3402 = write[1] ? n2378 : n1322;   // regs.v(46)
    assign n3403 = write[1] ? n2379 : n1323;   // regs.v(46)
    assign n3404 = write[1] ? n2380 : n1324;   // regs.v(46)
    assign n3405 = write[1] ? n2381 : n1325;   // regs.v(46)
    assign n3406 = write[1] ? n2382 : n1326;   // regs.v(46)
    assign n3407 = write[1] ? n2383 : n1327;   // regs.v(46)
    assign n3408 = write[1] ? n2384 : n1328;   // regs.v(46)
    assign n3409 = write[1] ? n2385 : n1329;   // regs.v(46)
    assign n3410 = write[1] ? n2386 : n1330;   // regs.v(46)
    assign n3411 = write[1] ? n2387 : n1331;   // regs.v(46)
    assign n3412 = write[1] ? n2388 : n1332;   // regs.v(46)
    assign n3413 = write[1] ? n2389 : n1333;   // regs.v(46)
    assign n3414 = write[1] ? n2390 : n1334;   // regs.v(46)
    assign n3415 = write[1] ? n2391 : n1335;   // regs.v(46)
    assign n3416 = write[1] ? n2392 : n1336;   // regs.v(46)
    assign n3417 = write[1] ? n2393 : n1337;   // regs.v(46)
    assign n3418 = write[1] ? n2394 : n1338;   // regs.v(46)
    assign n3419 = write[1] ? n2395 : n1339;   // regs.v(46)
    assign n3420 = write[1] ? n2396 : n1340;   // regs.v(46)
    assign n3421 = write[1] ? n2397 : n1341;   // regs.v(46)
    assign n3422 = write[1] ? n2398 : n1342;   // regs.v(46)
    assign n3423 = write[1] ? n2399 : n1343;   // regs.v(46)
    assign n3424 = write[1] ? n2400 : n1344;   // regs.v(46)
    assign n3425 = write[1] ? n2401 : n1345;   // regs.v(46)
    assign n3426 = write[1] ? n2402 : n1346;   // regs.v(46)
    assign n3427 = write[1] ? n2403 : n1347;   // regs.v(46)
    assign n3428 = write[1] ? n2404 : n1348;   // regs.v(46)
    assign n3429 = write[1] ? n2405 : n1349;   // regs.v(46)
    assign n3430 = write[1] ? n2406 : n1350;   // regs.v(46)
    assign n3431 = write[1] ? n2407 : n1351;   // regs.v(46)
    assign n3432 = write[1] ? n2408 : n1352;   // regs.v(46)
    assign n3433 = write[1] ? n2409 : n1353;   // regs.v(46)
    assign n3434 = write[1] ? n2410 : n1354;   // regs.v(46)
    assign n3435 = write[1] ? n2411 : n1355;   // regs.v(46)
    assign n3436 = write[1] ? n2412 : n1356;   // regs.v(46)
    assign n3437 = write[1] ? n2413 : n1357;   // regs.v(46)
    assign n3438 = write[1] ? n2414 : n1358;   // regs.v(46)
    assign n3439 = write[1] ? n2415 : n1359;   // regs.v(46)
    assign n3440 = write[1] ? n2416 : n1360;   // regs.v(46)
    assign n3441 = write[1] ? n2417 : n1361;   // regs.v(46)
    assign n3442 = write[1] ? n2418 : n1362;   // regs.v(46)
    assign n3443 = write[1] ? n2419 : n1363;   // regs.v(46)
    assign n3444 = write[1] ? n2420 : n1364;   // regs.v(46)
    assign n3445 = write[1] ? n2421 : n1365;   // regs.v(46)
    assign n3446 = write[1] ? n2422 : n1366;   // regs.v(46)
    assign n3447 = write[1] ? n2423 : n1367;   // regs.v(46)
    assign n3448 = write[1] ? n2424 : n1368;   // regs.v(46)
    assign n3449 = write[1] ? n2425 : n1369;   // regs.v(46)
    assign n3450 = write[1] ? n2426 : n1370;   // regs.v(46)
    assign n3451 = write[1] ? n2427 : n1371;   // regs.v(46)
    assign n3452 = write[1] ? n2428 : n1372;   // regs.v(46)
    assign n3453 = write[1] ? n2429 : n1373;   // regs.v(46)
    assign n3454 = write[1] ? n2430 : n1374;   // regs.v(46)
    assign n3455 = write[1] ? n2431 : n1375;   // regs.v(46)
    assign n3456 = write[1] ? n2432 : n1376;   // regs.v(46)
    assign n3457 = write[1] ? n2433 : n1377;   // regs.v(46)
    assign n3458 = write[1] ? n2434 : n1378;   // regs.v(46)
    assign n3459 = write[1] ? n2435 : n1379;   // regs.v(46)
    assign n3460 = write[1] ? n2436 : n1380;   // regs.v(46)
    assign n3461 = write[1] ? n2437 : n1381;   // regs.v(46)
    assign n3462 = write[1] ? n2438 : n1382;   // regs.v(46)
    assign n3463 = write[1] ? n2439 : n1383;   // regs.v(46)
    assign n3464 = write[1] ? n2440 : n1384;   // regs.v(46)
    assign n3465 = write[1] ? n2441 : n1385;   // regs.v(46)
    assign n3466 = write[1] ? n2442 : n1386;   // regs.v(46)
    assign n3467 = write[1] ? n2443 : n1387;   // regs.v(46)
    assign n3468 = write[1] ? n2444 : n1388;   // regs.v(46)
    assign n3469 = write[1] ? n2445 : n1389;   // regs.v(46)
    assign n3470 = write[1] ? n2446 : n1390;   // regs.v(46)
    assign n3471 = write[1] ? n2447 : n1391;   // regs.v(46)
    assign n3472 = write[1] ? n2448 : n1392;   // regs.v(46)
    assign n3473 = write[1] ? n2449 : n1393;   // regs.v(46)
    assign n3474 = write[1] ? n2450 : n1394;   // regs.v(46)
    assign n3475 = write[1] ? n2451 : n1395;   // regs.v(46)
    assign n3476 = write[1] ? n2452 : n1396;   // regs.v(46)
    assign n3477 = write[1] ? n2453 : n1397;   // regs.v(46)
    assign n3478 = write[1] ? n2454 : n1398;   // regs.v(46)
    assign n3479 = write[1] ? n2455 : n1399;   // regs.v(46)
    assign n3480 = write[1] ? n2456 : n1400;   // regs.v(46)
    assign n3481 = write[1] ? n2457 : n1401;   // regs.v(46)
    assign n3482 = write[1] ? n2458 : n1402;   // regs.v(46)
    assign n3483 = write[1] ? n2459 : n1403;   // regs.v(46)
    assign n3484 = write[1] ? n2460 : n1404;   // regs.v(46)
    assign n3485 = write[1] ? n2461 : n1405;   // regs.v(46)
    assign n3486 = write[1] ? n2462 : n1406;   // regs.v(46)
    assign n3487 = write[1] ? n2463 : n1407;   // regs.v(46)
    assign n3488 = write[1] ? n2464 : n1408;   // regs.v(46)
    assign n3489 = write[1] ? n2465 : n1409;   // regs.v(46)
    assign n3490 = write[1] ? n2466 : n1410;   // regs.v(46)
    assign n3491 = write[1] ? n2467 : n1411;   // regs.v(46)
    assign n3492 = write[1] ? n2468 : n1412;   // regs.v(46)
    assign n3493 = write[1] ? n2469 : n1413;   // regs.v(46)
    assign n3494 = write[1] ? n2470 : n1414;   // regs.v(46)
    assign n3495 = write[1] ? n2471 : n1415;   // regs.v(46)
    assign n3496 = write[1] ? n2472 : n1416;   // regs.v(46)
    assign n3497 = write[1] ? n2473 : n1417;   // regs.v(46)
    assign n3498 = write[1] ? n2474 : n1418;   // regs.v(46)
    assign n3499 = write[1] ? n2475 : n1419;   // regs.v(46)
    assign n3500 = write[1] ? n2476 : n1420;   // regs.v(46)
    assign n3501 = write[1] ? n2477 : n1421;   // regs.v(46)
    assign n3502 = write[1] ? n2478 : n1422;   // regs.v(46)
    assign n3503 = write[1] ? n2479 : n1423;   // regs.v(46)
    assign n3504 = write[1] ? n2480 : n1424;   // regs.v(46)
    assign n3505 = write[1] ? n2481 : n1425;   // regs.v(46)
    assign n3506 = write[1] ? n2482 : n1426;   // regs.v(46)
    assign n3507 = write[1] ? n2483 : n1427;   // regs.v(46)
    assign n3508 = write[1] ? n2484 : n1428;   // regs.v(46)
    assign n3509 = write[1] ? n2485 : n1429;   // regs.v(46)
    assign n3510 = write[1] ? n2486 : n1430;   // regs.v(46)
    assign n3511 = write[1] ? n2487 : n1431;   // regs.v(46)
    assign n3512 = write[1] ? n2488 : n1432;   // regs.v(46)
    assign n3513 = write[1] ? n2489 : n1433;   // regs.v(46)
    assign n3514 = write[1] ? n2490 : n1434;   // regs.v(46)
    assign n3515 = write[1] ? n2491 : n1435;   // regs.v(46)
    assign n3516 = write[1] ? n2492 : n1436;   // regs.v(46)
    assign n3517 = write[1] ? n2493 : n1437;   // regs.v(46)
    assign n3518 = write[1] ? n2494 : n1438;   // regs.v(46)
    assign n3519 = write[1] ? n2495 : n1439;   // regs.v(46)
    assign n3520 = write[1] ? n2496 : n1440;   // regs.v(46)
    assign n3521 = write[1] ? n2497 : n1441;   // regs.v(46)
    assign n3522 = write[1] ? n2498 : n1442;   // regs.v(46)
    assign n3523 = write[1] ? n2499 : n1443;   // regs.v(46)
    assign n3524 = write[1] ? n2500 : n1444;   // regs.v(46)
    assign n3525 = write[1] ? n2501 : n1445;   // regs.v(46)
    assign n3526 = write[1] ? n2502 : n1446;   // regs.v(46)
    assign n3527 = write[1] ? n2503 : n1447;   // regs.v(46)
    assign n3528 = write[1] ? n2504 : n1448;   // regs.v(46)
    assign n3529 = write[1] ? n2505 : n1449;   // regs.v(46)
    assign n3530 = write[1] ? n2506 : n1450;   // regs.v(46)
    assign n3531 = write[1] ? n2507 : n1451;   // regs.v(46)
    assign n3532 = write[1] ? n2508 : n1452;   // regs.v(46)
    assign n3533 = write[1] ? n2509 : n1453;   // regs.v(46)
    assign n3534 = write[1] ? n2510 : n1454;   // regs.v(46)
    assign n3535 = write[1] ? n2511 : n1455;   // regs.v(46)
    assign n3536 = write[1] ? n2512 : n1456;   // regs.v(46)
    assign n3537 = write[1] ? n2513 : n1457;   // regs.v(46)
    assign n3538 = write[1] ? n2514 : n1458;   // regs.v(46)
    assign n3539 = write[1] ? n2515 : n1459;   // regs.v(46)
    assign n3540 = write[1] ? n2516 : n1460;   // regs.v(46)
    assign n3541 = write[1] ? n2517 : n1461;   // regs.v(46)
    assign n3542 = write[1] ? n2518 : n1462;   // regs.v(46)
    assign n3543 = write[1] ? n2519 : n1463;   // regs.v(46)
    assign n3544 = write[1] ? n2520 : n1464;   // regs.v(46)
    assign n3545 = write[1] ? n2521 : n1465;   // regs.v(46)
    assign n3546 = write[1] ? n2522 : n1466;   // regs.v(46)
    assign n3547 = write[1] ? n2523 : n1467;   // regs.v(46)
    assign n3548 = write[1] ? n2524 : n1468;   // regs.v(46)
    assign n3549 = write[1] ? n2525 : n1469;   // regs.v(46)
    assign n3550 = write[1] ? n2526 : n1470;   // regs.v(46)
    assign n3551 = write[1] ? n2527 : n1471;   // regs.v(46)
    assign n3552 = write[1] ? n2528 : n1472;   // regs.v(46)
    assign n3553 = write[1] ? n2529 : n1473;   // regs.v(46)
    assign n3554 = write[1] ? n2530 : n1474;   // regs.v(46)
    assign n3555 = write[1] ? n2531 : n1475;   // regs.v(46)
    assign n3556 = write[1] ? n2532 : n1476;   // regs.v(46)
    assign n3557 = write[1] ? n2533 : n1477;   // regs.v(46)
    assign n3558 = write[1] ? n2534 : n1478;   // regs.v(46)
    assign n3559 = write[1] ? n2535 : n1479;   // regs.v(46)
    assign n3560 = write[1] ? n2536 : n1480;   // regs.v(46)
    assign n3561 = write[1] ? n2537 : n1481;   // regs.v(46)
    assign n3562 = write[1] ? n2538 : n1482;   // regs.v(46)
    assign n3563 = write[1] ? n2539 : n1483;   // regs.v(46)
    assign n3564 = write[1] ? n2540 : n1484;   // regs.v(46)
    assign n3565 = write[1] ? n2541 : n1485;   // regs.v(46)
    assign n3566 = write[1] ? n2542 : n1486;   // regs.v(46)
    assign n3567 = write[1] ? n2543 : n1487;   // regs.v(46)
    assign n3568 = write[1] ? n2544 : n1488;   // regs.v(46)
    assign n3569 = write[1] ? n2545 : n1489;   // regs.v(46)
    assign n3570 = write[1] ? n2546 : n1490;   // regs.v(46)
    assign n3571 = write[1] ? n2547 : n1491;   // regs.v(46)
    assign n3572 = write[1] ? n2548 : n1492;   // regs.v(46)
    assign n3573 = write[1] ? n2549 : n1493;   // regs.v(46)
    assign n3574 = write[1] ? n2550 : n1494;   // regs.v(46)
    assign n3575 = write[1] ? n2551 : n1495;   // regs.v(46)
    assign n3576 = write[1] ? n2552 : n1496;   // regs.v(46)
    assign n3577 = write[1] ? n2553 : n1497;   // regs.v(46)
    assign n3578 = write[1] ? n2554 : n1498;   // regs.v(46)
    assign n3579 = write[1] ? n2555 : n1499;   // regs.v(46)
    assign n3580 = write[1] ? n2556 : n1500;   // regs.v(46)
    assign n3581 = write[1] ? n2557 : n1501;   // regs.v(46)
    assign n3582 = write[1] ? n2558 : n1502;   // regs.v(46)
    assign n3583 = write[1] ? n2559 : n1503;   // regs.v(46)
    assign n3584 = write[1] ? n2560 : n1504;   // regs.v(46)
    assign n3585 = write[1] ? n2561 : n1505;   // regs.v(46)
    assign n3586 = write[1] ? n2562 : n1506;   // regs.v(46)
    assign n3587 = write[1] ? n2563 : n1507;   // regs.v(46)
    assign n3588 = write[1] ? n2564 : n1508;   // regs.v(46)
    assign n3589 = write[1] ? n2565 : n1509;   // regs.v(46)
    assign n3590 = write[1] ? n2566 : n1510;   // regs.v(46)
    assign n3591 = write[1] ? n2567 : n1511;   // regs.v(46)
    assign n3592 = write[1] ? n2568 : n1512;   // regs.v(46)
    assign n3593 = write[1] ? n2569 : n1513;   // regs.v(46)
    assign n3594 = write[1] ? n2570 : n1514;   // regs.v(46)
    assign n3595 = write[1] ? n2571 : n1515;   // regs.v(46)
    assign n3596 = write[1] ? n2572 : n1516;   // regs.v(46)
    assign n3597 = write[1] ? n2573 : n1517;   // regs.v(46)
    assign n3598 = write[1] ? n2574 : n1518;   // regs.v(46)
    assign n3599 = write[1] ? n2575 : n1519;   // regs.v(46)
    assign n3600 = write[1] ? n2576 : n1520;   // regs.v(46)
    assign n3601 = write[1] ? n2577 : n1521;   // regs.v(46)
    assign n3602 = write[1] ? n2578 : n1522;   // regs.v(46)
    assign n3603 = write[1] ? n2579 : n1523;   // regs.v(46)
    assign n3604 = write[1] ? n2580 : n1524;   // regs.v(46)
    assign n3605 = write[1] ? n2581 : n1525;   // regs.v(46)
    assign n3606 = write[1] ? n2582 : n1526;   // regs.v(46)
    assign n3607 = write[1] ? n2583 : n1527;   // regs.v(46)
    assign n3608 = write[1] ? n2584 : n1528;   // regs.v(46)
    assign n3609 = write[1] ? n2585 : n1529;   // regs.v(46)
    assign n3610 = write[1] ? n2586 : n1530;   // regs.v(46)
    assign n3611 = write[1] ? n2587 : n1531;   // regs.v(46)
    assign n3612 = write[1] ? n2588 : n1532;   // regs.v(46)
    assign n3613 = write[1] ? n2589 : n1533;   // regs.v(46)
    assign n3614 = write[1] ? n2590 : n1534;   // regs.v(46)
    assign n3615 = write[1] ? n2591 : n1535;   // regs.v(46)
    assign n3616 = write[1] ? n2592 : n1536;   // regs.v(46)
    assign n3617 = write[1] ? n2593 : n1537;   // regs.v(46)
    assign n3618 = write[1] ? n2594 : n1538;   // regs.v(46)
    assign n3619 = write[1] ? n2595 : n1539;   // regs.v(46)
    assign n3620 = write[1] ? n2596 : n1540;   // regs.v(46)
    assign n3621 = write[1] ? n2597 : n1541;   // regs.v(46)
    assign n3622 = write[1] ? n2598 : n1542;   // regs.v(46)
    assign n3623 = write[1] ? n2599 : n1543;   // regs.v(46)
    assign n3624 = write[1] ? n2600 : n1544;   // regs.v(46)
    assign n3625 = write[1] ? n2601 : n1545;   // regs.v(46)
    assign n3626 = write[1] ? n2602 : n1546;   // regs.v(46)
    assign n3627 = write[1] ? n2603 : n1547;   // regs.v(46)
    assign n3628 = write[1] ? n2604 : n1548;   // regs.v(46)
    assign n3629 = write[1] ? n2605 : n1549;   // regs.v(46)
    assign n3630 = write[1] ? n2606 : n1550;   // regs.v(46)
    assign n3631 = write[1] ? n2607 : n1551;   // regs.v(46)
    assign n3632 = write[1] ? n2608 : n1552;   // regs.v(46)
    assign n3633 = write[1] ? n2609 : n1553;   // regs.v(46)
    assign n3634 = write[1] ? n2610 : n1554;   // regs.v(46)
    assign n3635 = write[1] ? n2611 : n1555;   // regs.v(46)
    assign n3636 = write[1] ? n2612 : n1556;   // regs.v(46)
    assign n3637 = write[1] ? n2613 : n1557;   // regs.v(46)
    assign n3638 = write[1] ? n2614 : n1558;   // regs.v(46)
    assign n3639 = write[1] ? n2615 : n1559;   // regs.v(46)
    assign n3640 = write[1] ? n2616 : n1560;   // regs.v(46)
    assign n3641 = write[1] ? n2617 : n1561;   // regs.v(46)
    assign n3642 = write[1] ? n2618 : n1562;   // regs.v(46)
    assign n3643 = write[1] ? n2619 : n1563;   // regs.v(46)
    assign n3644 = write[1] ? n2620 : n1564;   // regs.v(46)
    assign n3645 = write[1] ? n2621 : n1565;   // regs.v(46)
    assign n3646 = write[1] ? n2622 : n1566;   // regs.v(46)
    assign n3647 = write[1] ? n2623 : n1567;   // regs.v(46)
    assign n3648 = write[1] ? n2624 : n1568;   // regs.v(46)
    assign n3649 = write[1] ? n2625 : n1569;   // regs.v(46)
    assign n3650 = write[1] ? n2626 : n1570;   // regs.v(46)
    assign n3651 = write[1] ? n2627 : n1571;   // regs.v(46)
    assign n3652 = write[1] ? n2628 : n1572;   // regs.v(46)
    assign n3653 = write[1] ? n2629 : n1573;   // regs.v(46)
    assign n3654 = write[1] ? n2630 : n1574;   // regs.v(46)
    assign n3655 = write[1] ? n2631 : n1575;   // regs.v(46)
    assign n3656 = write[1] ? n2632 : n1576;   // regs.v(46)
    assign n3657 = write[1] ? n2633 : n1577;   // regs.v(46)
    assign n3658 = write[1] ? n2634 : n1578;   // regs.v(46)
    assign n3659 = write[1] ? n2635 : n1579;   // regs.v(46)
    assign n3660 = write[1] ? n2636 : n1580;   // regs.v(46)
    assign n3661 = write[1] ? n2637 : n1581;   // regs.v(46)
    assign n3662 = write[1] ? n2638 : n1582;   // regs.v(46)
    assign n3663 = write[1] ? n2639 : n1583;   // regs.v(46)
    assign n3664 = write[1] ? n2640 : n1584;   // regs.v(46)
    assign n3665 = write[1] ? n2641 : n1585;   // regs.v(46)
    assign n3666 = write[1] ? n2642 : n1586;   // regs.v(46)
    assign n3667 = write[1] ? n2643 : n1587;   // regs.v(46)
    assign n3668 = write[1] ? n2644 : n1588;   // regs.v(46)
    assign n3669 = write[1] ? n2645 : n1589;   // regs.v(46)
    assign n3670 = write[1] ? n2646 : n1590;   // regs.v(46)
    assign n3671 = write[1] ? n2647 : n1591;   // regs.v(46)
    assign n3672 = write[1] ? n2648 : n1592;   // regs.v(46)
    assign n3673 = write[1] ? n2649 : n1593;   // regs.v(46)
    assign n3674 = write[1] ? n2650 : n1594;   // regs.v(46)
    assign n3675 = write[1] ? n2651 : n1595;   // regs.v(46)
    assign n3676 = write[1] ? n2652 : n1596;   // regs.v(46)
    assign n3677 = write[1] ? n2653 : n1597;   // regs.v(46)
    assign n3678 = write[1] ? n2654 : n1598;   // regs.v(46)
    assign n3679 = write[1] ? n2655 : n1599;   // regs.v(46)
    assign n3680 = write[1] ? n2656 : n1600;   // regs.v(46)
    assign n3681 = write[1] ? n2657 : n1601;   // regs.v(46)
    assign n3682 = write[1] ? n2658 : n1602;   // regs.v(46)
    assign n3683 = write[1] ? n2659 : n1603;   // regs.v(46)
    assign n3684 = write[1] ? n2660 : n1604;   // regs.v(46)
    assign n3685 = write[1] ? n2661 : n1605;   // regs.v(46)
    assign n3686 = write[1] ? n2662 : n1606;   // regs.v(46)
    assign n3687 = write[1] ? n2663 : n1607;   // regs.v(46)
    assign n3688 = write[1] ? n2664 : n1608;   // regs.v(46)
    assign n3689 = write[1] ? n2665 : n1609;   // regs.v(46)
    assign n3690 = write[1] ? n2666 : n1610;   // regs.v(46)
    assign n3691 = write[1] ? n2667 : n1611;   // regs.v(46)
    assign n3692 = write[1] ? n2668 : n1612;   // regs.v(46)
    assign n3693 = write[1] ? n2669 : n1613;   // regs.v(46)
    assign n3694 = write[1] ? n2670 : n1614;   // regs.v(46)
    assign n3695 = write[1] ? n2671 : n1615;   // regs.v(46)
    assign n3696 = write[1] ? n2672 : n1616;   // regs.v(46)
    assign n3697 = write[1] ? n2673 : n1617;   // regs.v(46)
    assign n3698 = write[1] ? n2674 : n1618;   // regs.v(46)
    assign n3699 = write[1] ? n2675 : n1619;   // regs.v(46)
    assign n3700 = write[1] ? n2676 : n1620;   // regs.v(46)
    assign n3701 = write[1] ? n2677 : n1621;   // regs.v(46)
    assign n3702 = write[1] ? n2678 : n1622;   // regs.v(46)
    assign n3703 = write[1] ? n2679 : n1623;   // regs.v(46)
    assign n3704 = write[1] ? n2680 : n1624;   // regs.v(46)
    assign n3705 = write[1] ? n2681 : n1625;   // regs.v(46)
    assign n3706 = write[1] ? n2682 : n1626;   // regs.v(46)
    assign n3707 = write[1] ? n2683 : n1627;   // regs.v(46)
    assign n3708 = write[1] ? n2684 : n1628;   // regs.v(46)
    assign n3709 = write[1] ? n2685 : n1629;   // regs.v(46)
    assign n3710 = write[1] ? n2686 : n1630;   // regs.v(46)
    assign n3711 = write[1] ? n2687 : n1631;   // regs.v(46)
    assign n3712 = write[1] ? n2688 : n1632;   // regs.v(46)
    assign n3713 = write[1] ? n2689 : n1633;   // regs.v(46)
    assign n3714 = write[1] ? n2690 : n1634;   // regs.v(46)
    assign n3715 = write[1] ? n2691 : n1635;   // regs.v(46)
    assign n3716 = write[1] ? n2692 : n1636;   // regs.v(46)
    assign n3717 = write[1] ? n2693 : n1637;   // regs.v(46)
    assign n3718 = write[1] ? n2694 : n1638;   // regs.v(46)
    assign n3719 = write[1] ? n2695 : n1639;   // regs.v(46)
    assign n3720 = write[1] ? n2696 : n1640;   // regs.v(46)
    assign n3721 = write[1] ? n2697 : n1641;   // regs.v(46)
    assign n3722 = write[1] ? n2698 : n1642;   // regs.v(46)
    assign n3723 = write[1] ? n2699 : n1643;   // regs.v(46)
    assign n3724 = write[1] ? n2700 : n1644;   // regs.v(46)
    assign n3725 = write[1] ? n2701 : n1645;   // regs.v(46)
    assign n3726 = write[1] ? n2702 : n1646;   // regs.v(46)
    assign n3727 = write[1] ? n2703 : n1647;   // regs.v(46)
    assign n3728 = write[1] ? n2704 : n1648;   // regs.v(46)
    assign n3729 = write[1] ? n2705 : n1649;   // regs.v(46)
    assign n3730 = write[1] ? n2706 : n1650;   // regs.v(46)
    assign n3731 = write[1] ? n2707 : n1651;   // regs.v(46)
    assign n3732 = write[1] ? n2708 : n1652;   // regs.v(46)
    assign n3733 = write[1] ? n2709 : n1653;   // regs.v(46)
    assign n3734 = write[1] ? n2710 : n1654;   // regs.v(46)
    assign n3735 = write[1] ? n2711 : n1655;   // regs.v(46)
    assign n3736 = write[1] ? n2712 : n1656;   // regs.v(46)
    assign n3737 = write[1] ? n2713 : n1657;   // regs.v(46)
    assign n3738 = write[1] ? n2714 : n1658;   // regs.v(46)
    assign n3739 = write[1] ? n2715 : n1659;   // regs.v(46)
    assign n3740 = write[1] ? n2716 : n1660;   // regs.v(46)
    assign n3741 = write[1] ? n2717 : n1661;   // regs.v(46)
    assign n3742 = write[1] ? n2718 : n1662;   // regs.v(46)
    assign n3743 = write[1] ? n2719 : n1663;   // regs.v(46)
    assign n3744 = write[1] ? n2720 : n1664;   // regs.v(46)
    assign n3745 = write[1] ? n2721 : n1665;   // regs.v(46)
    assign n3746 = write[1] ? n2722 : n1666;   // regs.v(46)
    assign n3747 = write[1] ? n2723 : n1667;   // regs.v(46)
    assign n3748 = write[1] ? n2724 : n1668;   // regs.v(46)
    assign n3749 = write[1] ? n2725 : n1669;   // regs.v(46)
    assign n3750 = write[1] ? n2726 : n1670;   // regs.v(46)
    assign n3751 = write[1] ? n2727 : n1671;   // regs.v(46)
    assign n3752 = write[1] ? n2728 : n1672;   // regs.v(46)
    assign n3753 = write[1] ? n2729 : n1673;   // regs.v(46)
    assign n3754 = write[1] ? n2730 : n1674;   // regs.v(46)
    assign n3755 = write[1] ? n2731 : n1675;   // regs.v(46)
    assign n3756 = write[1] ? n2732 : n1676;   // regs.v(46)
    assign n3757 = write[1] ? n2733 : n1677;   // regs.v(46)
    assign n3758 = write[1] ? n2734 : n1678;   // regs.v(46)
    assign n3759 = write[1] ? n2735 : n1679;   // regs.v(46)
    assign n3760 = write[1] ? n2736 : n1680;   // regs.v(46)
    assign n3761 = write[1] ? n2737 : n1681;   // regs.v(46)
    assign n3762 = write[1] ? n2738 : n1682;   // regs.v(46)
    assign n3763 = write[1] ? n2739 : n1683;   // regs.v(46)
    assign n3764 = write[1] ? n2740 : n1684;   // regs.v(46)
    assign n3765 = write[1] ? n2741 : n1685;   // regs.v(46)
    assign n3766 = write[1] ? n2742 : n1686;   // regs.v(46)
    assign n3767 = write[1] ? n2743 : n1687;   // regs.v(46)
    assign n3768 = write[1] ? n2744 : n1688;   // regs.v(46)
    assign n3769 = write[1] ? n2745 : n1689;   // regs.v(46)
    assign n3770 = write[1] ? n2746 : n1690;   // regs.v(46)
    assign n3771 = write[1] ? n2747 : n1691;   // regs.v(46)
    assign n3772 = write[1] ? n2748 : n1692;   // regs.v(46)
    assign n3773 = write[1] ? n2749 : n1693;   // regs.v(46)
    assign n3774 = write[1] ? n2750 : n1694;   // regs.v(46)
    assign n3775 = write[1] ? n2751 : n1695;   // regs.v(46)
    assign n3776 = write[1] ? n2752 : n1696;   // regs.v(46)
    assign n3777 = write[1] ? n2753 : n1697;   // regs.v(46)
    assign n3778 = write[1] ? n2754 : n1698;   // regs.v(46)
    assign n3779 = write[1] ? n2755 : n1699;   // regs.v(46)
    assign n3780 = write[1] ? n2756 : n1700;   // regs.v(46)
    assign n3781 = write[1] ? n2757 : n1701;   // regs.v(46)
    assign n3782 = write[1] ? n2758 : n1702;   // regs.v(46)
    assign n3783 = write[1] ? n2759 : n1703;   // regs.v(46)
    assign n3784 = write[1] ? n2760 : n1704;   // regs.v(46)
    assign n3785 = write[1] ? n2761 : n1705;   // regs.v(46)
    assign n3786 = write[1] ? n2762 : n1706;   // regs.v(46)
    assign n3787 = write[1] ? n2763 : n1707;   // regs.v(46)
    assign n3788 = write[1] ? n2764 : n1708;   // regs.v(46)
    assign n3789 = write[1] ? n2765 : n1709;   // regs.v(46)
    assign n3790 = write[1] ? n2766 : n1710;   // regs.v(46)
    assign n3791 = write[1] ? n2767 : n1711;   // regs.v(46)
    assign n3792 = write[1] ? n2768 : n1712;   // regs.v(46)
    assign n3793 = write[1] ? n2769 : n1713;   // regs.v(46)
    assign n3794 = write[1] ? n2770 : n1714;   // regs.v(46)
    assign n3795 = write[1] ? n2771 : n1715;   // regs.v(46)
    assign n3796 = write[1] ? n2772 : n1716;   // regs.v(46)
    assign n3797 = write[1] ? n2773 : n1717;   // regs.v(46)
    assign n3798 = write[1] ? n2774 : n1718;   // regs.v(46)
    assign n3799 = write[1] ? n2775 : n1719;   // regs.v(46)
    assign n3800 = write[1] ? n2776 : n1720;   // regs.v(46)
    assign n3801 = write[1] ? n2777 : n1721;   // regs.v(46)
    assign n3802 = write[1] ? n2778 : n1722;   // regs.v(46)
    assign n3803 = write[1] ? n2779 : n1723;   // regs.v(46)
    assign n3804 = write[1] ? n2780 : n1724;   // regs.v(46)
    assign n3805 = write[1] ? n2781 : n1725;   // regs.v(46)
    assign n3806 = write[1] ? n2782 : n1726;   // regs.v(46)
    assign n3807 = write[1] ? n2783 : n1727;   // regs.v(46)
    assign n3808 = write[1] ? n2784 : n1728;   // regs.v(46)
    assign n3809 = write[1] ? n2785 : n1729;   // regs.v(46)
    assign n3810 = write[1] ? n2786 : n1730;   // regs.v(46)
    assign n3811 = write[1] ? n2787 : n1731;   // regs.v(46)
    assign n3812 = write[1] ? n2788 : n1732;   // regs.v(46)
    assign n3813 = write[1] ? n2789 : n1733;   // regs.v(46)
    assign n3814 = write[1] ? n2790 : n1734;   // regs.v(46)
    assign n3815 = write[1] ? n2791 : n1735;   // regs.v(46)
    assign n3816 = write[1] ? n2792 : n1736;   // regs.v(46)
    assign n3817 = write[1] ? n2793 : n1737;   // regs.v(46)
    assign n3818 = write[1] ? n2794 : n1738;   // regs.v(46)
    assign n3819 = write[1] ? n2795 : n1739;   // regs.v(46)
    assign n3820 = write[1] ? n2796 : n1740;   // regs.v(46)
    assign n3821 = write[1] ? n2797 : n1741;   // regs.v(46)
    assign n3822 = write[1] ? n2798 : n1742;   // regs.v(46)
    assign n3823 = write[1] ? n2799 : n1743;   // regs.v(46)
    assign n3824 = write[1] ? n2800 : n1744;   // regs.v(46)
    assign n3825 = write[1] ? n2801 : n1745;   // regs.v(46)
    assign n3826 = write[1] ? n2802 : n1746;   // regs.v(46)
    assign n3827 = write[1] ? n2803 : n1747;   // regs.v(46)
    assign n3828 = write[1] ? n2804 : n1748;   // regs.v(46)
    assign n3829 = write[1] ? n2805 : n1749;   // regs.v(46)
    assign n3830 = write[1] ? n2806 : n1750;   // regs.v(46)
    assign n3831 = write[1] ? n2807 : n1751;   // regs.v(46)
    assign n3832 = write[1] ? n2808 : n1752;   // regs.v(46)
    assign n3833 = write[1] ? n2809 : n1753;   // regs.v(46)
    assign n3834 = write[1] ? n2810 : n1754;   // regs.v(46)
    assign n3835 = write[1] ? n2811 : n1755;   // regs.v(46)
    assign n3836 = write[1] ? n2812 : n1756;   // regs.v(46)
    assign n3837 = write[1] ? n2813 : n1757;   // regs.v(46)
    assign n3838 = write[1] ? n2814 : n1758;   // regs.v(46)
    assign n3839 = write[1] ? n2815 : n1759;   // regs.v(46)
    assign n3840 = write[1] ? n2816 : n1760;   // regs.v(46)
    assign n3841 = write[1] ? n2817 : n1761;   // regs.v(46)
    assign n3842 = write[1] ? n2818 : n1762;   // regs.v(46)
    assign n3843 = write[1] ? n2819 : n1763;   // regs.v(46)
    assign n3844 = write[1] ? n2820 : n1764;   // regs.v(46)
    assign n3845 = write[1] ? n2821 : n1765;   // regs.v(46)
    assign n3846 = write[1] ? n2822 : n1766;   // regs.v(46)
    assign n3847 = write[1] ? n2823 : n1767;   // regs.v(46)
    assign n3848 = write[1] ? n2824 : n1768;   // regs.v(46)
    assign n3849 = write[1] ? n2825 : n1769;   // regs.v(46)
    assign n3850 = write[1] ? n2826 : n1770;   // regs.v(46)
    assign n3851 = write[1] ? n2827 : n1771;   // regs.v(46)
    assign n3852 = write[1] ? n2828 : n1772;   // regs.v(46)
    assign n3853 = write[1] ? n2829 : n1773;   // regs.v(46)
    assign n3854 = write[1] ? n2830 : n1774;   // regs.v(46)
    assign n3855 = write[1] ? n2831 : n1775;   // regs.v(46)
    assign n3856 = write[1] ? n2832 : n1776;   // regs.v(46)
    assign n3857 = write[1] ? n2833 : n1777;   // regs.v(46)
    assign n3858 = write[1] ? n2834 : n1778;   // regs.v(46)
    assign n3859 = write[1] ? n2835 : n1779;   // regs.v(46)
    assign n3860 = write[1] ? n2836 : n1780;   // regs.v(46)
    assign n3861 = write[1] ? n2837 : n1781;   // regs.v(46)
    assign n3862 = write[1] ? n2838 : n1782;   // regs.v(46)
    assign n3863 = write[1] ? n2839 : n1783;   // regs.v(46)
    assign n3864 = write[1] ? n2840 : n1784;   // regs.v(46)
    assign n3865 = write[1] ? n2841 : n1785;   // regs.v(46)
    assign n3866 = write[1] ? n2842 : n1786;   // regs.v(46)
    assign n3867 = write[1] ? n2843 : n1787;   // regs.v(46)
    assign n3868 = write[1] ? n2844 : n1788;   // regs.v(46)
    assign n3869 = write[1] ? n2845 : n1789;   // regs.v(46)
    assign n3870 = write[1] ? n2846 : n1790;   // regs.v(46)
    assign n3871 = write[1] ? n2847 : n1791;   // regs.v(46)
    assign n3872 = write[1] ? n2848 : n1792;   // regs.v(46)
    assign n3873 = write[1] ? n2849 : n1793;   // regs.v(46)
    assign n3874 = write[1] ? n2850 : n1794;   // regs.v(46)
    assign n3875 = write[1] ? n2851 : n1795;   // regs.v(46)
    assign n3876 = write[1] ? n2852 : n1796;   // regs.v(46)
    assign n3877 = write[1] ? n2853 : n1797;   // regs.v(46)
    assign n3878 = write[1] ? n2854 : n1798;   // regs.v(46)
    assign n3879 = write[1] ? n2855 : n1799;   // regs.v(46)
    assign n3880 = write[1] ? n2856 : n1800;   // regs.v(46)
    assign n3881 = write[1] ? n2857 : n1801;   // regs.v(46)
    assign n3882 = write[1] ? n2858 : n1802;   // regs.v(46)
    assign n3883 = write[1] ? n2859 : n1803;   // regs.v(46)
    assign n3884 = write[1] ? n2860 : n1804;   // regs.v(46)
    assign n3885 = write[1] ? n2861 : n1805;   // regs.v(46)
    assign n3886 = write[1] ? n2862 : n1806;   // regs.v(46)
    assign n3887 = write[1] ? n2863 : n1807;   // regs.v(46)
    assign n3888 = write[1] ? n2864 : n1808;   // regs.v(46)
    assign n3889 = write[1] ? n2865 : n1809;   // regs.v(46)
    assign n3890 = write[1] ? n2866 : n1810;   // regs.v(46)
    assign n3891 = write[1] ? n2867 : n1811;   // regs.v(46)
    assign n3892 = write[1] ? n2868 : n1812;   // regs.v(46)
    assign n3893 = write[1] ? n2869 : n1813;   // regs.v(46)
    assign n3894 = write[1] ? n2870 : n1814;   // regs.v(46)
    assign n3895 = write[1] ? n2871 : n1815;   // regs.v(46)
    assign n3896 = write[1] ? n2872 : n1816;   // regs.v(46)
    assign n3897 = write[1] ? n2873 : n1817;   // regs.v(46)
    assign n3898 = write[1] ? n2874 : n1818;   // regs.v(46)
    assign n3899 = write[1] ? n2875 : n1819;   // regs.v(46)
    assign n3900 = write[1] ? n2876 : n1820;   // regs.v(46)
    assign n3901 = write[1] ? n2877 : n1821;   // regs.v(46)
    assign n3902 = write[1] ? n2878 : n1822;   // regs.v(46)
    assign n3903 = write[1] ? n2879 : n1823;   // regs.v(46)
    assign n3904 = write[1] ? n2880 : n1824;   // regs.v(46)
    assign n3905 = write[1] ? n2881 : n1825;   // regs.v(46)
    assign n3906 = write[1] ? n2882 : n1826;   // regs.v(46)
    assign n3907 = write[1] ? n2883 : n1827;   // regs.v(46)
    assign n3908 = write[1] ? n2884 : n1828;   // regs.v(46)
    assign n3909 = write[1] ? n2885 : n1829;   // regs.v(46)
    assign n3910 = write[1] ? n2886 : n1830;   // regs.v(46)
    assign n3911 = write[1] ? n2887 : n1831;   // regs.v(46)
    assign n3912 = write[1] ? n2888 : n1832;   // regs.v(46)
    assign n3913 = write[1] ? n2889 : n1833;   // regs.v(46)
    assign n3914 = write[1] ? n2890 : n1834;   // regs.v(46)
    assign n3915 = write[1] ? n2891 : n1835;   // regs.v(46)
    assign n3916 = write[1] ? n2892 : n1836;   // regs.v(46)
    assign n3917 = write[1] ? n2893 : n1837;   // regs.v(46)
    assign n3918 = write[1] ? n2894 : n1838;   // regs.v(46)
    assign n3919 = write[1] ? n2895 : n1839;   // regs.v(46)
    assign n3920 = write[1] ? n2896 : n1840;   // regs.v(46)
    assign n3921 = write[1] ? n2897 : n1841;   // regs.v(46)
    assign n3922 = write[1] ? n2898 : n1842;   // regs.v(46)
    assign n3923 = write[1] ? n2899 : n1843;   // regs.v(46)
    assign n3924 = write[1] ? n2900 : n1844;   // regs.v(46)
    assign n3925 = write[1] ? n2901 : n1845;   // regs.v(46)
    assign n3926 = write[1] ? n2902 : n1846;   // regs.v(46)
    assign n3927 = write[1] ? n2903 : n1847;   // regs.v(46)
    assign n3928 = write[1] ? n2904 : n1848;   // regs.v(46)
    assign n3929 = write[1] ? n2905 : n1849;   // regs.v(46)
    assign n3930 = write[1] ? n2906 : n1850;   // regs.v(46)
    assign n3931 = write[1] ? n2907 : n1851;   // regs.v(46)
    assign n3932 = write[1] ? n2908 : n1852;   // regs.v(46)
    assign n3933 = write[1] ? n2909 : n1853;   // regs.v(46)
    assign n3934 = write[1] ? n2910 : n1854;   // regs.v(46)
    assign n3935 = write[1] ? n2911 : n1855;   // regs.v(46)
    assign n3936 = write[1] ? n2912 : n1856;   // regs.v(46)
    assign n3937 = write[1] ? n2913 : n1857;   // regs.v(46)
    assign n3938 = write[1] ? n2914 : n1858;   // regs.v(46)
    assign n3939 = write[1] ? n2915 : n1859;   // regs.v(46)
    assign n3940 = write[1] ? n2916 : n1860;   // regs.v(46)
    assign n3941 = write[1] ? n2917 : n1861;   // regs.v(46)
    assign n3942 = write[1] ? n2918 : n1862;   // regs.v(46)
    assign n3943 = write[1] ? n2919 : n1863;   // regs.v(46)
    assign n3944 = write[1] ? n2920 : n1864;   // regs.v(46)
    assign n3945 = write[1] ? n2921 : n1865;   // regs.v(46)
    assign n3946 = write[1] ? n2922 : n1866;   // regs.v(46)
    assign n3947 = write[1] ? n2923 : n1867;   // regs.v(46)
    assign n3948 = write[1] ? n2924 : n1868;   // regs.v(46)
    assign n3949 = write[1] ? n2925 : n1869;   // regs.v(46)
    assign n3950 = write[1] ? n2926 : n1870;   // regs.v(46)
    assign n3951 = write[1] ? n2927 : n1871;   // regs.v(46)
    assign n3952 = write[1] ? n2928 : n1872;   // regs.v(46)
    assign n3953 = write[1] ? n2929 : n1873;   // regs.v(46)
    assign n3954 = write[1] ? n2930 : n1874;   // regs.v(46)
    assign n3955 = write[1] ? n2931 : n1875;   // regs.v(46)
    assign n3956 = write[1] ? n2932 : n1876;   // regs.v(46)
    assign n3957 = write[1] ? n2933 : n1877;   // regs.v(46)
    assign n3958 = write[1] ? n2934 : n1878;   // regs.v(46)
    assign n3959 = write[1] ? n2935 : n1879;   // regs.v(46)
    assign n3960 = write[1] ? n2936 : n1880;   // regs.v(46)
    assign n3961 = write[1] ? n2937 : n1881;   // regs.v(46)
    assign n3962 = write[1] ? n2938 : n1882;   // regs.v(46)
    assign n3963 = write[1] ? n2939 : n1883;   // regs.v(46)
    assign n3964 = write[1] ? n2940 : n1884;   // regs.v(46)
    assign n3965 = write[1] ? n2941 : n1885;   // regs.v(46)
    assign n3966 = write[1] ? n2942 : n1886;   // regs.v(46)
    assign n3967 = write[1] ? n2943 : n1887;   // regs.v(46)
    assign n3968 = write[1] ? n2944 : n1888;   // regs.v(46)
    assign n3969 = write[1] ? n2945 : n1889;   // regs.v(46)
    assign n3970 = write[1] ? n2946 : n1890;   // regs.v(46)
    assign n3971 = write[1] ? n2947 : n1891;   // regs.v(46)
    assign n3972 = write[1] ? n2948 : n1892;   // regs.v(46)
    assign n3973 = write[1] ? n2949 : n1893;   // regs.v(46)
    assign n3974 = write[1] ? n2950 : n1894;   // regs.v(46)
    assign n3975 = write[1] ? n2951 : n1895;   // regs.v(46)
    assign n3976 = write[1] ? n2952 : n1896;   // regs.v(46)
    assign n3977 = write[1] ? n2953 : n1897;   // regs.v(46)
    assign n3978 = write[1] ? n2954 : n1898;   // regs.v(46)
    assign n3979 = write[1] ? n2955 : n1899;   // regs.v(46)
    assign n3980 = write[1] ? n2956 : n1900;   // regs.v(46)
    assign n3981 = write[1] ? n2957 : n1901;   // regs.v(46)
    assign n3982 = write[1] ? n2958 : n1902;   // regs.v(46)
    assign n3983 = write[1] ? n2959 : n1903;   // regs.v(46)
    assign n3984 = write[1] ? n2960 : n1904;   // regs.v(46)
    assign n3985 = write[1] ? n2961 : n1905;   // regs.v(46)
    assign n3986 = write[1] ? n2962 : n1906;   // regs.v(46)
    assign n3987 = write[1] ? n2963 : n1907;   // regs.v(46)
    assign n3988 = write[1] ? n2964 : n1908;   // regs.v(46)
    assign n3989 = write[1] ? n2965 : n1909;   // regs.v(46)
    assign n3990 = write[1] ? n2966 : n1910;   // regs.v(46)
    assign n3991 = write[1] ? n2967 : n1911;   // regs.v(46)
    assign n3992 = write[1] ? n2968 : n1912;   // regs.v(46)
    assign n3993 = write[1] ? n2969 : n1913;   // regs.v(46)
    assign n3994 = write[1] ? n2970 : n1914;   // regs.v(46)
    assign n3995 = write[1] ? n2971 : n1915;   // regs.v(46)
    assign n3996 = write[1] ? n2972 : n1916;   // regs.v(46)
    assign n3997 = write[1] ? n2973 : n1917;   // regs.v(46)
    assign n3998 = write[1] ? n2974 : n1918;   // regs.v(46)
    assign n3999 = write[1] ? n2975 : n1919;   // regs.v(46)
    assign n4000 = write[1] ? n2976 : n1920;   // regs.v(46)
    assign n4001 = write[1] ? n2977 : n1921;   // regs.v(46)
    assign n4002 = write[1] ? n2978 : n1922;   // regs.v(46)
    assign n4003 = write[1] ? n2979 : n1923;   // regs.v(46)
    assign n4004 = write[1] ? n2980 : n1924;   // regs.v(46)
    assign n4005 = write[1] ? n2981 : n1925;   // regs.v(46)
    assign n4006 = write[1] ? n2982 : n1926;   // regs.v(46)
    assign n4007 = write[1] ? n2983 : n1927;   // regs.v(46)
    assign n4008 = write[1] ? n2984 : n1928;   // regs.v(46)
    assign n4009 = write[1] ? n2985 : n1929;   // regs.v(46)
    assign n4010 = write[1] ? n2986 : n1930;   // regs.v(46)
    assign n4011 = write[1] ? n2987 : n1931;   // regs.v(46)
    assign n4012 = write[1] ? n2988 : n1932;   // regs.v(46)
    assign n4013 = write[1] ? n2989 : n1933;   // regs.v(46)
    assign n4014 = write[1] ? n2990 : n1934;   // regs.v(46)
    assign n4015 = write[1] ? n2991 : n1935;   // regs.v(46)
    assign n4016 = write[1] ? n2992 : n1936;   // regs.v(46)
    assign n4017 = write[1] ? n2993 : n1937;   // regs.v(46)
    assign n4018 = write[1] ? n2994 : n1938;   // regs.v(46)
    assign n4019 = write[1] ? n2995 : n1939;   // regs.v(46)
    assign n4020 = write[1] ? n2996 : n1940;   // regs.v(46)
    assign n4021 = write[1] ? n2997 : n1941;   // regs.v(46)
    assign n4022 = write[1] ? n2998 : n1942;   // regs.v(46)
    assign n4023 = write[1] ? n2999 : n1943;   // regs.v(46)
    assign n4024 = write[1] ? n3000 : n1944;   // regs.v(46)
    assign n4025 = write[1] ? n3001 : n1945;   // regs.v(46)
    assign n4026 = write[1] ? n3002 : n1946;   // regs.v(46)
    assign n4027 = write[1] ? n3003 : n1947;   // regs.v(46)
    assign n4028 = write[1] ? n3004 : n1948;   // regs.v(46)
    assign n4029 = write[1] ? n3005 : n1949;   // regs.v(46)
    assign n4030 = write[1] ? n3006 : n1950;   // regs.v(46)
    assign n4031 = write[1] ? n3007 : n1951;   // regs.v(46)
    assign n4032 = write[1] ? n3008 : n1952;   // regs.v(46)
    assign n4033 = write[1] ? n3009 : n1953;   // regs.v(46)
    assign n4034 = write[1] ? n3010 : n1954;   // regs.v(46)
    assign n4035 = write[1] ? n3011 : n1955;   // regs.v(46)
    assign n4036 = write[1] ? n3012 : n1956;   // regs.v(46)
    assign n4037 = write[1] ? n3013 : n1957;   // regs.v(46)
    assign n4038 = write[1] ? n3014 : n1958;   // regs.v(46)
    assign n4039 = write[1] ? n3015 : n1959;   // regs.v(46)
    assign n4040 = write[1] ? n3016 : n1960;   // regs.v(46)
    assign n4041 = write[1] ? n3017 : n1961;   // regs.v(46)
    assign n4042 = write[1] ? n3018 : n1962;   // regs.v(46)
    assign n4043 = write[1] ? n3019 : n1963;   // regs.v(46)
    assign n4044 = write[1] ? n3020 : n1964;   // regs.v(46)
    assign n4045 = write[1] ? n3021 : n1965;   // regs.v(46)
    assign n4046 = write[1] ? n3022 : n1966;   // regs.v(46)
    assign n4047 = write[1] ? n3023 : n1967;   // regs.v(46)
    assign n4048 = write[1] ? n3024 : n1968;   // regs.v(46)
    assign n4049 = write[1] ? n3025 : n1969;   // regs.v(46)
    assign n4050 = write[1] ? n3026 : n1970;   // regs.v(46)
    assign n4051 = write[1] ? n3027 : n1971;   // regs.v(46)
    assign n4052 = write[1] ? n3028 : n1972;   // regs.v(46)
    assign n4053 = write[1] ? n3029 : n1973;   // regs.v(46)
    assign n4054 = write[1] ? n3030 : n1974;   // regs.v(46)
    assign n4055 = write[1] ? n3031 : n1975;   // regs.v(46)
    assign n4056 = write[1] ? n3032 : n1976;   // regs.v(46)
    assign n4057 = write[1] ? n3033 : n1977;   // regs.v(46)
    assign n4058 = write[1] ? n3034 : n1978;   // regs.v(46)
    assign n4059 = write[1] ? n3035 : n1979;   // regs.v(46)
    assign n4060 = write[1] ? n3036 : n1980;   // regs.v(46)
    assign n4061 = write[1] ? n3037 : n1981;   // regs.v(46)
    assign n4062 = write[1] ? n3038 : n1982;   // regs.v(46)
    assign n4063 = write[1] ? n3039 : n1983;   // regs.v(46)
    assign n4064 = write[1] ? n3040 : n1984;   // regs.v(46)
    assign n4065 = write[1] ? n3041 : n1985;   // regs.v(46)
    assign n4066 = write[1] ? n3042 : n1986;   // regs.v(46)
    assign n4067 = write[1] ? n3043 : n1987;   // regs.v(46)
    assign n4068 = write[1] ? n3044 : n1988;   // regs.v(46)
    assign n4069 = write[1] ? n3045 : n1989;   // regs.v(46)
    assign n4070 = write[1] ? n3046 : n1990;   // regs.v(46)
    assign n4071 = write[1] ? n3047 : n1991;   // regs.v(46)
    assign n4072 = write[1] ? n3048 : n1992;   // regs.v(46)
    assign n4073 = write[1] ? n3049 : n1993;   // regs.v(46)
    assign n4074 = write[1] ? n3050 : n1994;   // regs.v(46)
    assign n4075 = write[1] ? n3051 : n1995;   // regs.v(46)
    assign n4076 = write[1] ? n3052 : n1996;   // regs.v(46)
    assign n4077 = write[1] ? n3053 : n1997;   // regs.v(46)
    assign n4078 = write[1] ? n3054 : n1998;   // regs.v(46)
    assign n4079 = write[1] ? n3055 : n1999;   // regs.v(46)
    assign n4080 = write[1] ? n3056 : n2000;   // regs.v(46)
    assign n4081 = write[1] ? n3057 : n2001;   // regs.v(46)
    assign n4082 = write[1] ? n3058 : n2002;   // regs.v(46)
    assign n4083 = write[1] ? n3059 : n2003;   // regs.v(46)
    assign n4084 = write[1] ? n3060 : n2004;   // regs.v(46)
    assign n4085 = write[1] ? n3061 : n2005;   // regs.v(46)
    assign n4086 = write[1] ? n3062 : n2006;   // regs.v(46)
    assign n4087 = write[1] ? n3063 : n2007;   // regs.v(46)
    assign n4088 = write[1] ? n3064 : n2008;   // regs.v(46)
    assign n4089 = write[1] ? n3065 : n2009;   // regs.v(46)
    assign n4090 = write[1] ? n3066 : n2010;   // regs.v(46)
    assign n4091 = write[1] ? n3067 : n2011;   // regs.v(46)
    assign n4092 = write[1] ? n3068 : n2012;   // regs.v(46)
    assign n4093 = write[1] ? n3069 : n2013;   // regs.v(46)
    assign n4094 = write[1] ? n3070 : n2014;   // regs.v(46)
    assign n4095 = write[1] ? n3071 : n2015;   // regs.v(46)
    assign n4096 = write[1] ? n3072 : n2016;   // regs.v(46)
    assign n4097 = write[1] ? n3073 : n2017;   // regs.v(46)
    assign n4098 = write[1] ? n3074 : n2018;   // regs.v(46)
    assign n4099 = write[1] ? n3075 : n2019;   // regs.v(46)
    assign n4100 = write[1] ? n3076 : n2020;   // regs.v(46)
    assign n4101 = write[1] ? n3077 : n2021;   // regs.v(46)
    assign n4102 = write[1] ? n3078 : n2022;   // regs.v(46)
    assign n4103 = write[1] ? n3079 : n2023;   // regs.v(46)
    assign n4104 = write[1] ? n3080 : n2024;   // regs.v(46)
    assign n4105 = write[1] ? n3081 : n2025;   // regs.v(46)
    assign n4106 = write[1] ? n3082 : n2026;   // regs.v(46)
    assign n4107 = write[1] ? n3083 : n2027;   // regs.v(46)
    assign n4108 = write[1] ? n3084 : n2028;   // regs.v(46)
    assign n4109 = write[1] ? n3085 : n2029;   // regs.v(46)
    assign n4110 = write[1] ? n3086 : n2030;   // regs.v(46)
    assign n4111 = write[1] ? n3087 : n2031;   // regs.v(46)
    assign n4112 = write[1] ? n3088 : n2032;   // regs.v(46)
    assign n4113 = write[1] ? n3089 : n2033;   // regs.v(46)
    assign n4114 = write[1] ? n3090 : n2034;   // regs.v(46)
    assign n4115 = write[1] ? n3091 : n2035;   // regs.v(46)
    assign n4116 = write[1] ? n3092 : n2036;   // regs.v(46)
    assign n4117 = write[1] ? n3093 : n2037;   // regs.v(46)
    assign n4118 = write[1] ? n3094 : n2038;   // regs.v(46)
    assign n4119 = write[1] ? n3095 : n2039;   // regs.v(46)
    assign n4120 = write[1] ? n3096 : n2040;   // regs.v(46)
    assign n4121 = write[1] ? n3097 : n2041;   // regs.v(46)
    assign n4122 = write[1] ? n3098 : n2042;   // regs.v(46)
    assign n4123 = write[1] ? n3099 : n2043;   // regs.v(46)
    assign n4124 = write[1] ? n3100 : n2044;   // regs.v(46)
    assign n4125 = write[1] ? n3101 : n2045;   // regs.v(46)
    assign n4126 = write[1] ? n3102 : n2046;   // regs.v(46)
    assign n4127 = write[1] ? n3103 : n2047;   // regs.v(46)
    assign n4128 = write[1] ? n3104 : n2048;   // regs.v(46)
    assign n4129 = write[1] ? n3105 : n2049;   // regs.v(46)
    assign n4130 = write[1] ? n3106 : n2050;   // regs.v(46)
    assign n4131 = write[1] ? n3107 : n2051;   // regs.v(46)
    assign n4132 = write[1] ? n3108 : n2052;   // regs.v(46)
    assign n4133 = write[1] ? n3109 : n2053;   // regs.v(46)
    assign n4134 = write[1] ? n3110 : n2054;   // regs.v(46)
    assign n4135 = write[1] ? n3111 : n2055;   // regs.v(46)
    assign n4136 = write[1] ? n3112 : n2056;   // regs.v(46)
    assign n4137 = write[1] ? n3113 : n2057;   // regs.v(46)
    assign n4138 = write[1] ? n3114 : n2058;   // regs.v(46)
    assign n4139 = write[1] ? n3115 : n2059;   // regs.v(46)
    assign n4140 = write[1] ? n3116 : n2060;   // regs.v(46)
    assign n4141 = write[1] ? n3117 : n2061;   // regs.v(46)
    assign n4142 = write[1] ? n3118 : n2062;   // regs.v(46)
    assign n4143 = write[1] ? n3119 : n2063;   // regs.v(46)
    assign n4144 = write[1] ? n3120 : n2064;   // regs.v(46)
    assign n4145 = write[1] ? n3121 : n2065;   // regs.v(46)
    assign n4146 = write[1] ? n3122 : n2066;   // regs.v(46)
    assign n4147 = write[1] ? n3123 : n2067;   // regs.v(46)
    assign n4148 = write[1] ? n3124 : n2068;   // regs.v(46)
    assign n4149 = write[1] ? n3125 : n2069;   // regs.v(46)
    assign n4150 = write[1] ? n3126 : n2070;   // regs.v(46)
    assign n4151 = write[1] ? n3127 : n2071;   // regs.v(46)
    assign n4152 = write[1] ? n3128 : n2072;   // regs.v(46)
    assign n4153 = write[1] ? n3129 : n2073;   // regs.v(46)
    assign n4154 = write[1] ? n3130 : n2074;   // regs.v(46)
    assign n4155 = write[1] ? n3131 : n2075;   // regs.v(46)
    assign n4156 = write[1] ? n3132 : n2076;   // regs.v(46)
    assign n4157 = write[1] ? n3133 : n2077;   // regs.v(46)
    assign n4158 = write[1] ? n3134 : n2078;   // regs.v(46)
    assign n4159 = write[1] ? n3135 : n2079;   // regs.v(46)
    assign n4160 = write[1] ? n3136 : n2080;   // regs.v(46)
    assign n4161 = write[1] ? n3137 : n2081;   // regs.v(46)
    assign n4162 = write[1] ? n3138 : n2082;   // regs.v(46)
    assign n4163 = write[1] ? n3139 : n2083;   // regs.v(46)
    assign n4164 = write[1] ? n3140 : n2084;   // regs.v(46)
    assign n4165 = write[1] ? n3141 : n2085;   // regs.v(46)
    assign n4166 = write[1] ? n3142 : n2086;   // regs.v(46)
    assign n4167 = write[1] ? n3143 : n2087;   // regs.v(46)
    assign n4168 = write[1] ? n3144 : n2088;   // regs.v(46)
    assign n4169 = write[1] ? n3145 : n2089;   // regs.v(46)
    assign n4170 = write[1] ? n3146 : n2090;   // regs.v(46)
    assign n4171 = write[1] ? n3147 : n2091;   // regs.v(46)
    assign n4172 = write[1] ? n3148 : n2092;   // regs.v(46)
    assign n4173 = write[1] ? n3149 : n2093;   // regs.v(46)
    assign n4174 = write[1] ? n3150 : n2094;   // regs.v(46)
    assign n4175 = write[1] ? n3151 : n2095;   // regs.v(46)
    assign n4176 = write[1] ? n3152 : n2096;   // regs.v(46)
    assign n4177 = write[1] ? n3153 : n2097;   // regs.v(46)
    assign n4178 = write[1] ? n3154 : n2098;   // regs.v(46)
    assign n4179 = write[1] ? n3155 : n2099;   // regs.v(46)
    assign n4180 = write[1] ? n3156 : n2100;   // regs.v(46)
    assign n4181 = write[1] ? n3157 : n2101;   // regs.v(46)
    assign n4182 = write[1] ? n3158 : n2102;   // regs.v(46)
    assign n4183 = write[1] ? n3159 : n2103;   // regs.v(46)
    assign n4184 = write[1] ? n3160 : n2104;   // regs.v(46)
    assign n4185 = write[1] ? n3161 : n2105;   // regs.v(46)
    assign n4186 = write[1] ? n3162 : n2106;   // regs.v(46)
    assign n4187 = write[1] ? n3163 : n2107;   // regs.v(46)
    assign n4188 = write[1] ? n3164 : n2108;   // regs.v(46)
    assign n4189 = write[1] ? n3165 : n2109;   // regs.v(46)
    assign n4190 = write[1] ? n3166 : n2110;   // regs.v(46)
    assign n4191 = write[1] ? n3167 : n2111;   // regs.v(46)
    assign n4192 = write[1] ? n3168 : n2112;   // regs.v(46)
    assign n4193 = write[1] ? n3169 : n2113;   // regs.v(46)
    assign n4194 = write[1] ? n3170 : n2114;   // regs.v(46)
    assign n4195 = write[1] ? n3171 : n2115;   // regs.v(46)
    assign n4196 = write[1] ? n3172 : n2116;   // regs.v(46)
    assign n4197 = write[1] ? n3173 : n2117;   // regs.v(46)
    assign n4198 = write[1] ? n3174 : n2118;   // regs.v(46)
    assign n4199 = write[1] ? n3175 : n2119;   // regs.v(46)
    assign n4200 = write[1] ? n3176 : n2120;   // regs.v(46)
    assign n4201 = write[1] ? n3177 : n2121;   // regs.v(46)
    assign n4202 = write[1] ? n3178 : n2122;   // regs.v(46)
    assign n4203 = write[1] ? n3179 : n2123;   // regs.v(46)
    assign n4204 = write[1] ? n3180 : n2124;   // regs.v(46)
    assign n4205 = write[1] ? n3181 : n2125;   // regs.v(46)
    assign n4206 = write[1] ? n3182 : n2126;   // regs.v(46)
    assign n4207 = write[1] ? n3183 : n2127;   // regs.v(46)
    assign n4208 = write[1] ? n3184 : n2128;   // regs.v(46)
    assign n4209 = write[1] ? n3185 : n2129;   // regs.v(46)
    assign n4210 = write[1] ? n3186 : n2130;   // regs.v(46)
    assign n4211 = write[1] ? n3187 : n2131;   // regs.v(46)
    assign n4212 = write[1] ? n3188 : n2132;   // regs.v(46)
    assign n4213 = write[1] ? n3189 : n2133;   // regs.v(46)
    assign n4214 = write[1] ? n3190 : n2134;   // regs.v(46)
    assign n4215 = write[1] ? n3191 : n2135;   // regs.v(46)
    assign n4216 = write[1] ? n3192 : n2136;   // regs.v(46)
    assign n4217 = write[1] ? n3193 : n2137;   // regs.v(46)
    assign n4218 = write[1] ? n3194 : n2138;   // regs.v(46)
    assign n4219 = write[1] ? n3195 : n2139;   // regs.v(46)
    assign n4220 = write[1] ? n3196 : n2140;   // regs.v(46)
    assign n4221 = write[1] ? n3197 : n2141;   // regs.v(46)
    assign n4222 = write[1] ? n3198 : n2142;   // regs.v(46)
    assign n4223 = write[1] ? n3199 : n2143;   // regs.v(46)
    assign n4224 = write[1] ? n3200 : n2144;   // regs.v(46)
    assign n4225 = write[1] ? n3201 : n2145;   // regs.v(46)
    assign n4226 = write[1] ? n3202 : n2146;   // regs.v(46)
    assign n4227 = write[1] ? n3203 : n2147;   // regs.v(46)
    assign n4228 = write[1] ? n3204 : n2148;   // regs.v(46)
    assign n4229 = stwr ? stin[31] : n3301;   // regs.v(48)
    assign n4230 = stwr ? stin[30] : n3302;   // regs.v(48)
    assign n4231 = stwr ? stin[29] : n3303;   // regs.v(48)
    assign n4232 = stwr ? stin[28] : n3304;   // regs.v(48)
    assign n4233 = stwr ? stin[27] : n3305;   // regs.v(48)
    assign n4234 = stwr ? stin[26] : n3306;   // regs.v(48)
    assign n4235 = stwr ? stin[25] : n3307;   // regs.v(48)
    assign n4236 = stwr ? stin[24] : n3308;   // regs.v(48)
    assign n4237 = stwr ? stin[23] : n3309;   // regs.v(48)
    assign n4238 = stwr ? stin[22] : n3310;   // regs.v(48)
    assign n4239 = stwr ? stin[21] : n3311;   // regs.v(48)
    assign n4240 = stwr ? stin[20] : n3312;   // regs.v(48)
    assign n4241 = stwr ? stin[19] : n3313;   // regs.v(48)
    assign n4242 = stwr ? stin[18] : n3314;   // regs.v(48)
    assign n4243 = stwr ? stin[17] : n3315;   // regs.v(48)
    assign n4244 = stwr ? stin[16] : n3316;   // regs.v(48)
    assign n4245 = stwr ? stin[15] : n3317;   // regs.v(48)
    assign n4246 = stwr ? stin[14] : n3318;   // regs.v(48)
    assign n4247 = stwr ? stin[13] : n3319;   // regs.v(48)
    assign n4248 = stwr ? stin[12] : n3320;   // regs.v(48)
    assign n4249 = stwr ? stin[11] : n3321;   // regs.v(48)
    assign n4250 = stwr ? stin[10] : n3322;   // regs.v(48)
    assign n4251 = stwr ? stin[9] : n3323;   // regs.v(48)
    assign n4252 = stwr ? stin[8] : n3324;   // regs.v(48)
    assign n4253 = stwr ? stin[7] : n3325;   // regs.v(48)
    assign n4254 = stwr ? stin[6] : n3326;   // regs.v(48)
    assign n4255 = stwr ? stin[5] : n3327;   // regs.v(48)
    assign n4256 = stwr ? stin[4] : n3328;   // regs.v(48)
    assign n4257 = stwr ? stin[3] : n3329;   // regs.v(48)
    assign n4258 = stwr ? stin[2] : n3330;   // regs.v(48)
    assign n4259 = stwr ? stin[1] : n3331;   // regs.v(48)
    assign n4260 = stwr ? stin[0] : n3332;   // regs.v(48)
    add_32u_32u add_4198 (.cin(1'b0), .a({pcout}), .b({32'b00000000000000000000000000000001}), 
            .o({n4262, n4263, n4264, n4265, n4266, n4267, n4268, 
            n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, 
            n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, 
            n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, 
            n4293}));   // regs.v(49)
    assign n4294 = pcincr ? n4262 : n3205;   // regs.v(49)
    assign n4295 = pcincr ? n4263 : n3206;   // regs.v(49)
    assign n4296 = pcincr ? n4264 : n3207;   // regs.v(49)
    assign n4297 = pcincr ? n4265 : n3208;   // regs.v(49)
    assign n4298 = pcincr ? n4266 : n3209;   // regs.v(49)
    assign n4299 = pcincr ? n4267 : n3210;   // regs.v(49)
    assign n4300 = pcincr ? n4268 : n3211;   // regs.v(49)
    assign n4301 = pcincr ? n4269 : n3212;   // regs.v(49)
    assign n4302 = pcincr ? n4270 : n3213;   // regs.v(49)
    assign n4303 = pcincr ? n4271 : n3214;   // regs.v(49)
    assign n4304 = pcincr ? n4272 : n3215;   // regs.v(49)
    assign n4305 = pcincr ? n4273 : n3216;   // regs.v(49)
    assign n4306 = pcincr ? n4274 : n3217;   // regs.v(49)
    assign n4307 = pcincr ? n4275 : n3218;   // regs.v(49)
    assign n4308 = pcincr ? n4276 : n3219;   // regs.v(49)
    assign n4309 = pcincr ? n4277 : n3220;   // regs.v(49)
    assign n4310 = pcincr ? n4278 : n3221;   // regs.v(49)
    assign n4311 = pcincr ? n4279 : n3222;   // regs.v(49)
    assign n4312 = pcincr ? n4280 : n3223;   // regs.v(49)
    assign n4313 = pcincr ? n4281 : n3224;   // regs.v(49)
    assign n4314 = pcincr ? n4282 : n3225;   // regs.v(49)
    assign n4315 = pcincr ? n4283 : n3226;   // regs.v(49)
    assign n4316 = pcincr ? n4284 : n3227;   // regs.v(49)
    assign n4317 = pcincr ? n4285 : n3228;   // regs.v(49)
    assign n4318 = pcincr ? n4286 : n3229;   // regs.v(49)
    assign n4319 = pcincr ? n4287 : n3230;   // regs.v(49)
    assign n4320 = pcincr ? n4288 : n3231;   // regs.v(49)
    assign n4321 = pcincr ? n4289 : n3232;   // regs.v(49)
    assign n4322 = pcincr ? n4290 : n3233;   // regs.v(49)
    assign n4323 = pcincr ? n4291 : n3234;   // regs.v(49)
    assign n4324 = pcincr ? n4292 : n3235;   // regs.v(49)
    assign n4325 = pcincr ? n4293 : n3236;   // regs.v(49)
    VERIFIC_DFFRS i4233 (.d(n4295), .clk(clk), .s(1'b0), .r(rst), .q(pcout[30]));   // regs.v(41)
    VERIFIC_DFFRS i4234 (.d(n4296), .clk(clk), .s(1'b0), .r(rst), .q(pcout[29]));   // regs.v(41)
    VERIFIC_DFFRS i4235 (.d(n4297), .clk(clk), .s(1'b0), .r(rst), .q(pcout[28]));   // regs.v(41)
    VERIFIC_DFFRS i4236 (.d(n4298), .clk(clk), .s(1'b0), .r(rst), .q(pcout[27]));   // regs.v(41)
    VERIFIC_DFFRS i4237 (.d(n4299), .clk(clk), .s(1'b0), .r(rst), .q(pcout[26]));   // regs.v(41)
    VERIFIC_DFFRS i4238 (.d(n4300), .clk(clk), .s(1'b0), .r(rst), .q(pcout[25]));   // regs.v(41)
    VERIFIC_DFFRS i4239 (.d(n4301), .clk(clk), .s(1'b0), .r(rst), .q(pcout[24]));   // regs.v(41)
    VERIFIC_DFFRS i4240 (.d(n4302), .clk(clk), .s(1'b0), .r(rst), .q(pcout[23]));   // regs.v(41)
    VERIFIC_DFFRS i4241 (.d(n4303), .clk(clk), .s(1'b0), .r(rst), .q(pcout[22]));   // regs.v(41)
    VERIFIC_DFFRS i4242 (.d(n4304), .clk(clk), .s(1'b0), .r(rst), .q(pcout[21]));   // regs.v(41)
    VERIFIC_DFFRS i4243 (.d(n4305), .clk(clk), .s(1'b0), .r(rst), .q(pcout[20]));   // regs.v(41)
    VERIFIC_DFFRS i4244 (.d(n4306), .clk(clk), .s(1'b0), .r(rst), .q(pcout[19]));   // regs.v(41)
    VERIFIC_DFFRS i4245 (.d(n4307), .clk(clk), .s(1'b0), .r(rst), .q(pcout[18]));   // regs.v(41)
    VERIFIC_DFFRS i4246 (.d(n4308), .clk(clk), .s(1'b0), .r(rst), .q(pcout[17]));   // regs.v(41)
    VERIFIC_DFFRS i4247 (.d(n4309), .clk(clk), .s(1'b0), .r(rst), .q(pcout[16]));   // regs.v(41)
    VERIFIC_DFFRS i4248 (.d(n4310), .clk(clk), .s(1'b0), .r(rst), .q(pcout[15]));   // regs.v(41)
    VERIFIC_DFFRS i4249 (.d(n4311), .clk(clk), .s(1'b0), .r(rst), .q(pcout[14]));   // regs.v(41)
    VERIFIC_DFFRS i4250 (.d(n4312), .clk(clk), .s(1'b0), .r(rst), .q(pcout[13]));   // regs.v(41)
    VERIFIC_DFFRS i4251 (.d(n4313), .clk(clk), .s(1'b0), .r(rst), .q(pcout[12]));   // regs.v(41)
    VERIFIC_DFFRS i4252 (.d(n4314), .clk(clk), .s(1'b0), .r(rst), .q(pcout[11]));   // regs.v(41)
    VERIFIC_DFFRS i4253 (.d(n4315), .clk(clk), .s(1'b0), .r(rst), .q(pcout[10]));   // regs.v(41)
    VERIFIC_DFFRS i4254 (.d(n4316), .clk(clk), .s(1'b0), .r(rst), .q(pcout[9]));   // regs.v(41)
    VERIFIC_DFFRS i4255 (.d(n4317), .clk(clk), .s(1'b0), .r(rst), .q(pcout[8]));   // regs.v(41)
    VERIFIC_DFFRS i4256 (.d(n4318), .clk(clk), .s(1'b0), .r(rst), .q(pcout[7]));   // regs.v(41)
    VERIFIC_DFFRS i4257 (.d(n4319), .clk(clk), .s(1'b0), .r(rst), .q(pcout[6]));   // regs.v(41)
    VERIFIC_DFFRS i4258 (.d(n4320), .clk(clk), .s(1'b0), .r(rst), .q(pcout[5]));   // regs.v(41)
    VERIFIC_DFFRS i4259 (.d(n4321), .clk(clk), .s(1'b0), .r(rst), .q(pcout[4]));   // regs.v(41)
    VERIFIC_DFFRS i4260 (.d(n4322), .clk(clk), .s(1'b0), .r(rst), .q(pcout[3]));   // regs.v(41)
    VERIFIC_DFFRS i4261 (.d(n4323), .clk(clk), .s(1'b0), .r(rst), .q(pcout[2]));   // regs.v(41)
    VERIFIC_DFFRS i4262 (.d(n4324), .clk(clk), .s(1'b0), .r(rst), .q(pcout[1]));   // regs.v(41)
    VERIFIC_DFFRS i4263 (.d(n4325), .clk(clk), .s(1'b0), .r(rst), .q(pcout[0]));   // regs.v(41)
    VERIFIC_DFFRS i4264 (.d(n3237), .clk(clk), .s(1'b0), .r(rst), .q(spout[31]));   // regs.v(41)
    VERIFIC_DFFRS i4265 (.d(n3238), .clk(clk), .s(1'b0), .r(rst), .q(spout[30]));   // regs.v(41)
    VERIFIC_DFFRS i4266 (.d(n3239), .clk(clk), .s(1'b0), .r(rst), .q(spout[29]));   // regs.v(41)
    VERIFIC_DFFRS i4267 (.d(n3240), .clk(clk), .s(1'b0), .r(rst), .q(spout[28]));   // regs.v(41)
    VERIFIC_DFFRS i4268 (.d(n3241), .clk(clk), .s(1'b0), .r(rst), .q(spout[27]));   // regs.v(41)
    VERIFIC_DFFRS i4269 (.d(n3242), .clk(clk), .s(1'b0), .r(rst), .q(spout[26]));   // regs.v(41)
    VERIFIC_DFFRS i4270 (.d(n3243), .clk(clk), .s(1'b0), .r(rst), .q(spout[25]));   // regs.v(41)
    VERIFIC_DFFRS i4271 (.d(n3244), .clk(clk), .s(1'b0), .r(rst), .q(spout[24]));   // regs.v(41)
    VERIFIC_DFFRS i4272 (.d(n3245), .clk(clk), .s(1'b0), .r(rst), .q(spout[23]));   // regs.v(41)
    VERIFIC_DFFRS i4273 (.d(n3246), .clk(clk), .s(1'b0), .r(rst), .q(spout[22]));   // regs.v(41)
    VERIFIC_DFFRS i4274 (.d(n3247), .clk(clk), .s(1'b0), .r(rst), .q(spout[21]));   // regs.v(41)
    VERIFIC_DFFRS i4275 (.d(n3248), .clk(clk), .s(1'b0), .r(rst), .q(spout[20]));   // regs.v(41)
    VERIFIC_DFFRS i4276 (.d(n3249), .clk(clk), .s(1'b0), .r(rst), .q(spout[19]));   // regs.v(41)
    VERIFIC_DFFRS i4277 (.d(n3250), .clk(clk), .s(1'b0), .r(rst), .q(spout[18]));   // regs.v(41)
    VERIFIC_DFFRS i4278 (.d(n3251), .clk(clk), .s(1'b0), .r(rst), .q(spout[17]));   // regs.v(41)
    VERIFIC_DFFRS i4279 (.d(n3252), .clk(clk), .s(1'b0), .r(rst), .q(spout[16]));   // regs.v(41)
    VERIFIC_DFFRS i4280 (.d(n3253), .clk(clk), .s(1'b0), .r(rst), .q(spout[15]));   // regs.v(41)
    VERIFIC_DFFRS i4281 (.d(n3254), .clk(clk), .s(1'b0), .r(rst), .q(spout[14]));   // regs.v(41)
    VERIFIC_DFFRS i4282 (.d(n3255), .clk(clk), .s(1'b0), .r(rst), .q(spout[13]));   // regs.v(41)
    VERIFIC_DFFRS i4283 (.d(n3256), .clk(clk), .s(1'b0), .r(rst), .q(spout[12]));   // regs.v(41)
    VERIFIC_DFFRS i4284 (.d(n3257), .clk(clk), .s(1'b0), .r(rst), .q(spout[11]));   // regs.v(41)
    VERIFIC_DFFRS i4285 (.d(n3258), .clk(clk), .s(1'b0), .r(rst), .q(spout[10]));   // regs.v(41)
    VERIFIC_DFFRS i4286 (.d(n3259), .clk(clk), .s(1'b0), .r(rst), .q(spout[9]));   // regs.v(41)
    VERIFIC_DFFRS i4287 (.d(n3260), .clk(clk), .s(1'b0), .r(rst), .q(spout[8]));   // regs.v(41)
    VERIFIC_DFFRS i4288 (.d(n3261), .clk(clk), .s(1'b0), .r(rst), .q(spout[7]));   // regs.v(41)
    VERIFIC_DFFRS i4289 (.d(n3262), .clk(clk), .s(1'b0), .r(rst), .q(spout[6]));   // regs.v(41)
    VERIFIC_DFFRS i4290 (.d(n3263), .clk(clk), .s(1'b0), .r(rst), .q(spout[5]));   // regs.v(41)
    VERIFIC_DFFRS i4291 (.d(n3264), .clk(clk), .s(1'b0), .r(rst), .q(spout[4]));   // regs.v(41)
    VERIFIC_DFFRS i4292 (.d(n3265), .clk(clk), .s(1'b0), .r(rst), .q(spout[3]));   // regs.v(41)
    VERIFIC_DFFRS i4293 (.d(n3266), .clk(clk), .s(1'b0), .r(rst), .q(spout[2]));   // regs.v(41)
    VERIFIC_DFFRS i4294 (.d(n3267), .clk(clk), .s(1'b0), .r(rst), .q(spout[1]));   // regs.v(41)
    VERIFIC_DFFRS i4295 (.d(n3268), .clk(clk), .s(1'b0), .r(rst), .q(spout[0]));   // regs.v(41)
    VERIFIC_DFFRS i4296 (.d(n3269), .clk(clk), .s(1'b0), .r(rst), .q(lrout[31]));   // regs.v(41)
    VERIFIC_DFFRS i4297 (.d(n3270), .clk(clk), .s(1'b0), .r(rst), .q(lrout[30]));   // regs.v(41)
    VERIFIC_DFFRS i4298 (.d(n3271), .clk(clk), .s(1'b0), .r(rst), .q(lrout[29]));   // regs.v(41)
    VERIFIC_DFFRS i4299 (.d(n3272), .clk(clk), .s(1'b0), .r(rst), .q(lrout[28]));   // regs.v(41)
    VERIFIC_DFFRS i4300 (.d(n3273), .clk(clk), .s(1'b0), .r(rst), .q(lrout[27]));   // regs.v(41)
    VERIFIC_DFFRS i4301 (.d(n3274), .clk(clk), .s(1'b0), .r(rst), .q(lrout[26]));   // regs.v(41)
    VERIFIC_DFFRS i4302 (.d(n3275), .clk(clk), .s(1'b0), .r(rst), .q(lrout[25]));   // regs.v(41)
    VERIFIC_DFFRS i4303 (.d(n3276), .clk(clk), .s(1'b0), .r(rst), .q(lrout[24]));   // regs.v(41)
    VERIFIC_DFFRS i4304 (.d(n3277), .clk(clk), .s(1'b0), .r(rst), .q(lrout[23]));   // regs.v(41)
    VERIFIC_DFFRS i4305 (.d(n3278), .clk(clk), .s(1'b0), .r(rst), .q(lrout[22]));   // regs.v(41)
    VERIFIC_DFFRS i4306 (.d(n3279), .clk(clk), .s(1'b0), .r(rst), .q(lrout[21]));   // regs.v(41)
    VERIFIC_DFFRS i4307 (.d(n3280), .clk(clk), .s(1'b0), .r(rst), .q(lrout[20]));   // regs.v(41)
    VERIFIC_DFFRS i4308 (.d(n3281), .clk(clk), .s(1'b0), .r(rst), .q(lrout[19]));   // regs.v(41)
    VERIFIC_DFFRS i4309 (.d(n3282), .clk(clk), .s(1'b0), .r(rst), .q(lrout[18]));   // regs.v(41)
    VERIFIC_DFFRS i4310 (.d(n3283), .clk(clk), .s(1'b0), .r(rst), .q(lrout[17]));   // regs.v(41)
    VERIFIC_DFFRS i4311 (.d(n3284), .clk(clk), .s(1'b0), .r(rst), .q(lrout[16]));   // regs.v(41)
    VERIFIC_DFFRS i4312 (.d(n3285), .clk(clk), .s(1'b0), .r(rst), .q(lrout[15]));   // regs.v(41)
    VERIFIC_DFFRS i4313 (.d(n3286), .clk(clk), .s(1'b0), .r(rst), .q(lrout[14]));   // regs.v(41)
    VERIFIC_DFFRS i4314 (.d(n3287), .clk(clk), .s(1'b0), .r(rst), .q(lrout[13]));   // regs.v(41)
    VERIFIC_DFFRS i4315 (.d(n3288), .clk(clk), .s(1'b0), .r(rst), .q(lrout[12]));   // regs.v(41)
    VERIFIC_DFFRS i4316 (.d(n3289), .clk(clk), .s(1'b0), .r(rst), .q(lrout[11]));   // regs.v(41)
    VERIFIC_DFFRS i4317 (.d(n3290), .clk(clk), .s(1'b0), .r(rst), .q(lrout[10]));   // regs.v(41)
    VERIFIC_DFFRS i4318 (.d(n3291), .clk(clk), .s(1'b0), .r(rst), .q(lrout[9]));   // regs.v(41)
    VERIFIC_DFFRS i4319 (.d(n3292), .clk(clk), .s(1'b0), .r(rst), .q(lrout[8]));   // regs.v(41)
    VERIFIC_DFFRS i4320 (.d(n3293), .clk(clk), .s(1'b0), .r(rst), .q(lrout[7]));   // regs.v(41)
    VERIFIC_DFFRS i4321 (.d(n3294), .clk(clk), .s(1'b0), .r(rst), .q(lrout[6]));   // regs.v(41)
    VERIFIC_DFFRS i4322 (.d(n3295), .clk(clk), .s(1'b0), .r(rst), .q(lrout[5]));   // regs.v(41)
    VERIFIC_DFFRS i4323 (.d(n3296), .clk(clk), .s(1'b0), .r(rst), .q(lrout[4]));   // regs.v(41)
    VERIFIC_DFFRS i4324 (.d(n3297), .clk(clk), .s(1'b0), .r(rst), .q(lrout[3]));   // regs.v(41)
    VERIFIC_DFFRS i4325 (.d(n3298), .clk(clk), .s(1'b0), .r(rst), .q(lrout[2]));   // regs.v(41)
    VERIFIC_DFFRS i4326 (.d(n3299), .clk(clk), .s(1'b0), .r(rst), .q(lrout[1]));   // regs.v(41)
    VERIFIC_DFFRS i4327 (.d(n3300), .clk(clk), .s(1'b0), .r(rst), .q(lrout[0]));   // regs.v(41)
    VERIFIC_DFFRS i4328 (.d(n4229), .clk(clk), .s(1'b0), .r(rst), .q(stout[31]));   // regs.v(41)
    VERIFIC_DFFRS i4329 (.d(n4230), .clk(clk), .s(1'b0), .r(rst), .q(stout[30]));   // regs.v(41)
    VERIFIC_DFFRS i4330 (.d(n4231), .clk(clk), .s(1'b0), .r(rst), .q(stout[29]));   // regs.v(41)
    VERIFIC_DFFRS i4331 (.d(n4232), .clk(clk), .s(1'b0), .r(rst), .q(stout[28]));   // regs.v(41)
    VERIFIC_DFFRS i4332 (.d(n4233), .clk(clk), .s(1'b0), .r(rst), .q(stout[27]));   // regs.v(41)
    VERIFIC_DFFRS i4333 (.d(n4234), .clk(clk), .s(1'b0), .r(rst), .q(stout[26]));   // regs.v(41)
    VERIFIC_DFFRS i4334 (.d(n4235), .clk(clk), .s(1'b0), .r(rst), .q(stout[25]));   // regs.v(41)
    VERIFIC_DFFRS i4335 (.d(n4236), .clk(clk), .s(1'b0), .r(rst), .q(stout[24]));   // regs.v(41)
    VERIFIC_DFFRS i4336 (.d(n4237), .clk(clk), .s(1'b0), .r(rst), .q(stout[23]));   // regs.v(41)
    VERIFIC_DFFRS i4337 (.d(n4238), .clk(clk), .s(1'b0), .r(rst), .q(stout[22]));   // regs.v(41)
    VERIFIC_DFFRS i4338 (.d(n4239), .clk(clk), .s(1'b0), .r(rst), .q(stout[21]));   // regs.v(41)
    VERIFIC_DFFRS i4339 (.d(n4240), .clk(clk), .s(1'b0), .r(rst), .q(stout[20]));   // regs.v(41)
    VERIFIC_DFFRS i4340 (.d(n4241), .clk(clk), .s(1'b0), .r(rst), .q(stout[19]));   // regs.v(41)
    VERIFIC_DFFRS i4341 (.d(n4242), .clk(clk), .s(1'b0), .r(rst), .q(stout[18]));   // regs.v(41)
    VERIFIC_DFFRS i4342 (.d(n4243), .clk(clk), .s(1'b0), .r(rst), .q(stout[17]));   // regs.v(41)
    VERIFIC_DFFRS i4343 (.d(n4244), .clk(clk), .s(1'b0), .r(rst), .q(stout[16]));   // regs.v(41)
    VERIFIC_DFFRS i4344 (.d(n4245), .clk(clk), .s(1'b0), .r(rst), .q(stout[15]));   // regs.v(41)
    VERIFIC_DFFRS i4345 (.d(n4246), .clk(clk), .s(1'b0), .r(rst), .q(stout[14]));   // regs.v(41)
    VERIFIC_DFFRS i4346 (.d(n4247), .clk(clk), .s(1'b0), .r(rst), .q(stout[13]));   // regs.v(41)
    VERIFIC_DFFRS i4347 (.d(n4248), .clk(clk), .s(1'b0), .r(rst), .q(stout[12]));   // regs.v(41)
    VERIFIC_DFFRS i4348 (.d(n4249), .clk(clk), .s(1'b0), .r(rst), .q(stout[11]));   // regs.v(41)
    VERIFIC_DFFRS i4349 (.d(n4250), .clk(clk), .s(1'b0), .r(rst), .q(stout[10]));   // regs.v(41)
    VERIFIC_DFFRS i4350 (.d(n4251), .clk(clk), .s(1'b0), .r(rst), .q(stout[9]));   // regs.v(41)
    VERIFIC_DFFRS i4351 (.d(n4252), .clk(clk), .s(1'b0), .r(rst), .q(stout[8]));   // regs.v(41)
    VERIFIC_DFFRS i4352 (.d(n4253), .clk(clk), .s(1'b0), .r(rst), .q(stout[7]));   // regs.v(41)
    VERIFIC_DFFRS i4353 (.d(n4254), .clk(clk), .s(1'b0), .r(rst), .q(stout[6]));   // regs.v(41)
    VERIFIC_DFFRS i4354 (.d(n4255), .clk(clk), .s(1'b0), .r(rst), .q(stout[5]));   // regs.v(41)
    VERIFIC_DFFRS i4355 (.d(n4256), .clk(clk), .s(1'b0), .r(rst), .q(stout[4]));   // regs.v(41)
    VERIFIC_DFFRS i4356 (.d(n4257), .clk(clk), .s(1'b0), .r(rst), .q(stout[3]));   // regs.v(41)
    VERIFIC_DFFRS i4357 (.d(n4258), .clk(clk), .s(1'b0), .r(rst), .q(stout[2]));   // regs.v(41)
    VERIFIC_DFFRS i4358 (.d(n4259), .clk(clk), .s(1'b0), .r(rst), .q(stout[1]));   // regs.v(41)
    VERIFIC_DFFRS i4359 (.d(n4260), .clk(clk), .s(1'b0), .r(rst), .q(stout[0]));   // regs.v(41)
    VERIFIC_DFFRS i4360 (.d(n3333), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4361 (.d(n3334), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4362 (.d(n3335), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4363 (.d(n3336), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4364 (.d(n3337), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4365 (.d(n3338), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4366 (.d(n3339), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4367 (.d(n3340), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4368 (.d(n3341), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4369 (.d(n3342), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4370 (.d(n3343), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4371 (.d(n3344), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4372 (.d(n3345), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4373 (.d(n3346), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4374 (.d(n3347), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4375 (.d(n3348), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4376 (.d(n3349), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4377 (.d(n3350), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4378 (.d(n3351), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4379 (.d(n3352), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4380 (.d(n3353), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4381 (.d(n3354), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4382 (.d(n3355), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4383 (.d(n3356), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4384 (.d(n3357), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4385 (.d(n3358), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4386 (.d(n3359), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4387 (.d(n3360), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4388 (.d(n3361), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4389 (.d(n3362), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4390 (.d(n3363), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4391 (.d(n3364), .clk(clk), .s(1'b0), .r(rst), .q(\regs[27] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4392 (.d(n3365), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4393 (.d(n3366), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4394 (.d(n3367), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4395 (.d(n3368), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4396 (.d(n3369), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4397 (.d(n3370), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4398 (.d(n3371), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4399 (.d(n3372), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4400 (.d(n3373), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4401 (.d(n3374), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4402 (.d(n3375), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4403 (.d(n3376), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4404 (.d(n3377), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4405 (.d(n3378), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4406 (.d(n3379), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4407 (.d(n3380), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4408 (.d(n3381), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4409 (.d(n3382), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4410 (.d(n3383), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4411 (.d(n3384), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4412 (.d(n3385), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4413 (.d(n3386), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4414 (.d(n3387), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4415 (.d(n3388), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4416 (.d(n3389), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4417 (.d(n3390), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4418 (.d(n3391), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4419 (.d(n3392), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4420 (.d(n3393), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4421 (.d(n3394), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4422 (.d(n3395), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4423 (.d(n3396), .clk(clk), .s(1'b0), .r(rst), .q(\regs[26] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4424 (.d(n3397), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4425 (.d(n3398), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4426 (.d(n3399), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4427 (.d(n3400), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4428 (.d(n3401), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4429 (.d(n3402), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4430 (.d(n3403), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4431 (.d(n3404), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4432 (.d(n3405), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4433 (.d(n3406), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4434 (.d(n3407), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4435 (.d(n3408), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4436 (.d(n3409), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4437 (.d(n3410), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4438 (.d(n3411), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4439 (.d(n3412), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4440 (.d(n3413), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4441 (.d(n3414), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4442 (.d(n3415), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4443 (.d(n3416), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4444 (.d(n3417), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4445 (.d(n3418), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4446 (.d(n3419), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4447 (.d(n3420), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4448 (.d(n3421), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4449 (.d(n3422), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4450 (.d(n3423), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4451 (.d(n3424), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4452 (.d(n3425), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4453 (.d(n3426), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4454 (.d(n3427), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4455 (.d(n3428), .clk(clk), .s(1'b0), .r(rst), .q(\regs[25] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4456 (.d(n3429), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4457 (.d(n3430), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4458 (.d(n3431), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4459 (.d(n3432), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4460 (.d(n3433), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4461 (.d(n3434), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4462 (.d(n3435), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4463 (.d(n3436), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4464 (.d(n3437), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4465 (.d(n3438), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4466 (.d(n3439), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4467 (.d(n3440), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4468 (.d(n3441), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4469 (.d(n3442), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4470 (.d(n3443), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4471 (.d(n3444), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4472 (.d(n3445), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4473 (.d(n3446), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4474 (.d(n3447), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4475 (.d(n3448), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4476 (.d(n3449), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4477 (.d(n3450), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4478 (.d(n3451), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4479 (.d(n3452), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4480 (.d(n3453), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4481 (.d(n3454), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4482 (.d(n3455), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4483 (.d(n3456), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4484 (.d(n3457), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4485 (.d(n3458), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4486 (.d(n3459), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4487 (.d(n3460), .clk(clk), .s(1'b0), .r(rst), .q(\regs[24] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4488 (.d(n3461), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4489 (.d(n3462), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4490 (.d(n3463), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4491 (.d(n3464), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4492 (.d(n3465), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4493 (.d(n3466), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4494 (.d(n3467), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4495 (.d(n3468), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4496 (.d(n3469), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4497 (.d(n3470), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4498 (.d(n3471), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4499 (.d(n3472), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4500 (.d(n3473), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4501 (.d(n3474), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4502 (.d(n3475), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4503 (.d(n3476), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4504 (.d(n3477), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4505 (.d(n3478), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4506 (.d(n3479), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4507 (.d(n3480), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4508 (.d(n3481), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4509 (.d(n3482), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4510 (.d(n3483), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4511 (.d(n3484), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4512 (.d(n3485), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4513 (.d(n3486), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4514 (.d(n3487), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4515 (.d(n3488), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4516 (.d(n3489), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4517 (.d(n3490), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4518 (.d(n3491), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4519 (.d(n3492), .clk(clk), .s(1'b0), .r(rst), .q(\regs[23] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4520 (.d(n3493), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4521 (.d(n3494), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4522 (.d(n3495), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4523 (.d(n3496), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4524 (.d(n3497), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4525 (.d(n3498), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4526 (.d(n3499), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4527 (.d(n3500), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4528 (.d(n3501), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4529 (.d(n3502), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4530 (.d(n3503), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4531 (.d(n3504), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4532 (.d(n3505), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4533 (.d(n3506), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4534 (.d(n3507), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4535 (.d(n3508), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4536 (.d(n3509), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4537 (.d(n3510), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4538 (.d(n3511), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4539 (.d(n3512), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4540 (.d(n3513), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4541 (.d(n3514), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4542 (.d(n3515), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4543 (.d(n3516), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4544 (.d(n3517), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4545 (.d(n3518), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4546 (.d(n3519), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4547 (.d(n3520), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4548 (.d(n3521), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4549 (.d(n3522), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4550 (.d(n3523), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4551 (.d(n3524), .clk(clk), .s(1'b0), .r(rst), .q(\regs[22] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4552 (.d(n3525), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4553 (.d(n3526), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4554 (.d(n3527), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4555 (.d(n3528), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4556 (.d(n3529), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4557 (.d(n3530), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4558 (.d(n3531), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4559 (.d(n3532), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4560 (.d(n3533), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4561 (.d(n3534), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4562 (.d(n3535), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4563 (.d(n3536), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4564 (.d(n3537), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4565 (.d(n3538), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4566 (.d(n3539), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4567 (.d(n3540), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4568 (.d(n3541), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4569 (.d(n3542), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4570 (.d(n3543), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4571 (.d(n3544), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4572 (.d(n3545), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4573 (.d(n3546), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4574 (.d(n3547), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4575 (.d(n3548), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4576 (.d(n3549), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4577 (.d(n3550), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4578 (.d(n3551), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4579 (.d(n3552), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4580 (.d(n3553), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4581 (.d(n3554), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4582 (.d(n3555), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4583 (.d(n3556), .clk(clk), .s(1'b0), .r(rst), .q(\regs[21] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4584 (.d(n3557), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4585 (.d(n3558), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4586 (.d(n3559), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4587 (.d(n3560), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4588 (.d(n3561), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4589 (.d(n3562), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4590 (.d(n3563), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4591 (.d(n3564), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4592 (.d(n3565), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4593 (.d(n3566), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4594 (.d(n3567), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4595 (.d(n3568), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4596 (.d(n3569), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4597 (.d(n3570), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4598 (.d(n3571), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4599 (.d(n3572), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4600 (.d(n3573), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4601 (.d(n3574), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4602 (.d(n3575), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4603 (.d(n3576), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4604 (.d(n3577), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4605 (.d(n3578), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4606 (.d(n3579), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4607 (.d(n3580), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4608 (.d(n3581), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4609 (.d(n3582), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4610 (.d(n3583), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4611 (.d(n3584), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4612 (.d(n3585), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4613 (.d(n3586), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4614 (.d(n3587), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4615 (.d(n3588), .clk(clk), .s(1'b0), .r(rst), .q(\regs[20] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4616 (.d(n3589), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4617 (.d(n3590), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4618 (.d(n3591), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4619 (.d(n3592), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4620 (.d(n3593), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4621 (.d(n3594), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4622 (.d(n3595), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4623 (.d(n3596), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4624 (.d(n3597), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4625 (.d(n3598), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4626 (.d(n3599), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4627 (.d(n3600), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4628 (.d(n3601), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4629 (.d(n3602), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4630 (.d(n3603), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4631 (.d(n3604), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4632 (.d(n3605), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4633 (.d(n3606), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4634 (.d(n3607), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4635 (.d(n3608), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4636 (.d(n3609), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4637 (.d(n3610), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4638 (.d(n3611), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4639 (.d(n3612), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4640 (.d(n3613), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4641 (.d(n3614), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4642 (.d(n3615), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4643 (.d(n3616), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4644 (.d(n3617), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4645 (.d(n3618), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4646 (.d(n3619), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4647 (.d(n3620), .clk(clk), .s(1'b0), .r(rst), .q(\regs[19] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4648 (.d(n3621), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4649 (.d(n3622), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4650 (.d(n3623), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4651 (.d(n3624), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4652 (.d(n3625), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4653 (.d(n3626), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4654 (.d(n3627), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4655 (.d(n3628), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4656 (.d(n3629), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4657 (.d(n3630), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4658 (.d(n3631), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4659 (.d(n3632), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4660 (.d(n3633), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4661 (.d(n3634), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4662 (.d(n3635), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4663 (.d(n3636), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4664 (.d(n3637), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4665 (.d(n3638), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4666 (.d(n3639), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4667 (.d(n3640), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4668 (.d(n3641), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4669 (.d(n3642), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4670 (.d(n3643), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4671 (.d(n3644), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4672 (.d(n3645), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4673 (.d(n3646), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4674 (.d(n3647), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4675 (.d(n3648), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4676 (.d(n3649), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4677 (.d(n3650), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4678 (.d(n3651), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4679 (.d(n3652), .clk(clk), .s(1'b0), .r(rst), .q(\regs[18] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4680 (.d(n3653), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4681 (.d(n3654), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4682 (.d(n3655), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4683 (.d(n3656), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4684 (.d(n3657), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4685 (.d(n3658), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4686 (.d(n3659), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4687 (.d(n3660), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4688 (.d(n3661), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4689 (.d(n3662), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4690 (.d(n3663), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4691 (.d(n3664), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4692 (.d(n3665), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4693 (.d(n3666), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4694 (.d(n3667), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4695 (.d(n3668), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4696 (.d(n3669), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4697 (.d(n3670), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4698 (.d(n3671), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4699 (.d(n3672), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4700 (.d(n3673), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4701 (.d(n3674), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4702 (.d(n3675), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4703 (.d(n3676), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4704 (.d(n3677), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4705 (.d(n3678), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4706 (.d(n3679), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4707 (.d(n3680), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4708 (.d(n3681), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4709 (.d(n3682), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4710 (.d(n3683), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4711 (.d(n3684), .clk(clk), .s(1'b0), .r(rst), .q(\regs[17] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4712 (.d(n3685), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4713 (.d(n3686), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4714 (.d(n3687), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4715 (.d(n3688), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4716 (.d(n3689), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4717 (.d(n3690), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4718 (.d(n3691), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4719 (.d(n3692), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4720 (.d(n3693), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4721 (.d(n3694), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4722 (.d(n3695), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4723 (.d(n3696), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4724 (.d(n3697), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4725 (.d(n3698), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4726 (.d(n3699), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4727 (.d(n3700), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4728 (.d(n3701), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4729 (.d(n3702), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4730 (.d(n3703), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4731 (.d(n3704), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4732 (.d(n3705), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4733 (.d(n3706), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4734 (.d(n3707), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4735 (.d(n3708), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4736 (.d(n3709), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4737 (.d(n3710), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4738 (.d(n3711), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4739 (.d(n3712), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4740 (.d(n3713), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4741 (.d(n3714), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4742 (.d(n3715), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4743 (.d(n3716), .clk(clk), .s(1'b0), .r(rst), .q(\regs[16] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4744 (.d(n3717), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4745 (.d(n3718), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4746 (.d(n3719), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4747 (.d(n3720), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4748 (.d(n3721), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4749 (.d(n3722), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4750 (.d(n3723), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4751 (.d(n3724), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4752 (.d(n3725), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4753 (.d(n3726), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4754 (.d(n3727), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4755 (.d(n3728), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4756 (.d(n3729), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4757 (.d(n3730), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4758 (.d(n3731), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4759 (.d(n3732), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4760 (.d(n3733), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4761 (.d(n3734), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4762 (.d(n3735), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4763 (.d(n3736), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4764 (.d(n3737), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4765 (.d(n3738), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4766 (.d(n3739), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4767 (.d(n3740), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4768 (.d(n3741), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4769 (.d(n3742), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4770 (.d(n3743), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4771 (.d(n3744), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4772 (.d(n3745), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4773 (.d(n3746), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4774 (.d(n3747), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4775 (.d(n3748), .clk(clk), .s(1'b0), .r(rst), .q(\regs[15] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4776 (.d(n3749), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4777 (.d(n3750), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4778 (.d(n3751), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4779 (.d(n3752), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4780 (.d(n3753), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4781 (.d(n3754), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4782 (.d(n3755), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4783 (.d(n3756), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4784 (.d(n3757), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4785 (.d(n3758), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4786 (.d(n3759), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4787 (.d(n3760), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4788 (.d(n3761), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4789 (.d(n3762), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4790 (.d(n3763), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4791 (.d(n3764), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4792 (.d(n3765), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4793 (.d(n3766), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4794 (.d(n3767), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4795 (.d(n3768), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4796 (.d(n3769), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4797 (.d(n3770), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4798 (.d(n3771), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4799 (.d(n3772), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4800 (.d(n3773), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4801 (.d(n3774), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4802 (.d(n3775), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4803 (.d(n3776), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4804 (.d(n3777), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4805 (.d(n3778), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4806 (.d(n3779), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4807 (.d(n3780), .clk(clk), .s(1'b0), .r(rst), .q(\regs[14] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4808 (.d(n3781), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4809 (.d(n3782), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4810 (.d(n3783), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4811 (.d(n3784), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4812 (.d(n3785), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4813 (.d(n3786), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4814 (.d(n3787), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4815 (.d(n3788), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4816 (.d(n3789), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4817 (.d(n3790), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4818 (.d(n3791), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4819 (.d(n3792), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4820 (.d(n3793), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4821 (.d(n3794), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4822 (.d(n3795), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4823 (.d(n3796), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4824 (.d(n3797), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4825 (.d(n3798), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4826 (.d(n3799), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4827 (.d(n3800), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4828 (.d(n3801), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4829 (.d(n3802), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4830 (.d(n3803), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4831 (.d(n3804), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4832 (.d(n3805), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4833 (.d(n3806), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4834 (.d(n3807), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4835 (.d(n3808), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4836 (.d(n3809), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4837 (.d(n3810), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4838 (.d(n3811), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4839 (.d(n3812), .clk(clk), .s(1'b0), .r(rst), .q(\regs[13] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4840 (.d(n3813), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4841 (.d(n3814), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4842 (.d(n3815), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4843 (.d(n3816), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4844 (.d(n3817), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4845 (.d(n3818), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4846 (.d(n3819), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4847 (.d(n3820), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4848 (.d(n3821), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4849 (.d(n3822), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4850 (.d(n3823), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4851 (.d(n3824), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4852 (.d(n3825), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4853 (.d(n3826), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4854 (.d(n3827), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4855 (.d(n3828), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4856 (.d(n3829), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4857 (.d(n3830), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4858 (.d(n3831), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4859 (.d(n3832), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4860 (.d(n3833), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4861 (.d(n3834), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4862 (.d(n3835), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4863 (.d(n3836), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4864 (.d(n3837), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4865 (.d(n3838), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4866 (.d(n3839), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4867 (.d(n3840), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4868 (.d(n3841), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4869 (.d(n3842), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4870 (.d(n3843), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4871 (.d(n3844), .clk(clk), .s(1'b0), .r(rst), .q(\regs[12] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4872 (.d(n3845), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4873 (.d(n3846), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4874 (.d(n3847), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4875 (.d(n3848), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4876 (.d(n3849), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4877 (.d(n3850), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4878 (.d(n3851), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4879 (.d(n3852), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4880 (.d(n3853), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4881 (.d(n3854), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4882 (.d(n3855), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4883 (.d(n3856), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4884 (.d(n3857), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4885 (.d(n3858), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4886 (.d(n3859), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4887 (.d(n3860), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4888 (.d(n3861), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4889 (.d(n3862), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4890 (.d(n3863), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4891 (.d(n3864), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4892 (.d(n3865), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4893 (.d(n3866), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4894 (.d(n3867), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4895 (.d(n3868), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4896 (.d(n3869), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4897 (.d(n3870), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4898 (.d(n3871), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4899 (.d(n3872), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4900 (.d(n3873), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4901 (.d(n3874), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4902 (.d(n3875), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4903 (.d(n3876), .clk(clk), .s(1'b0), .r(rst), .q(\regs[11] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4904 (.d(n3877), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4905 (.d(n3878), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4906 (.d(n3879), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4907 (.d(n3880), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4908 (.d(n3881), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4909 (.d(n3882), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4910 (.d(n3883), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4911 (.d(n3884), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4912 (.d(n3885), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4913 (.d(n3886), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4914 (.d(n3887), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4915 (.d(n3888), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4916 (.d(n3889), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4917 (.d(n3890), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4918 (.d(n3891), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4919 (.d(n3892), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4920 (.d(n3893), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4921 (.d(n3894), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4922 (.d(n3895), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4923 (.d(n3896), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4924 (.d(n3897), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4925 (.d(n3898), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4926 (.d(n3899), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4927 (.d(n3900), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4928 (.d(n3901), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4929 (.d(n3902), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4930 (.d(n3903), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4931 (.d(n3904), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4932 (.d(n3905), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4933 (.d(n3906), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4934 (.d(n3907), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4935 (.d(n3908), .clk(clk), .s(1'b0), .r(rst), .q(\regs[10] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4936 (.d(n3909), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4937 (.d(n3910), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4938 (.d(n3911), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4939 (.d(n3912), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4940 (.d(n3913), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4941 (.d(n3914), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4942 (.d(n3915), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4943 (.d(n3916), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4944 (.d(n3917), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4945 (.d(n3918), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4946 (.d(n3919), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4947 (.d(n3920), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4948 (.d(n3921), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4949 (.d(n3922), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4950 (.d(n3923), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4951 (.d(n3924), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4952 (.d(n3925), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4953 (.d(n3926), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4954 (.d(n3927), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4955 (.d(n3928), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4956 (.d(n3929), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4957 (.d(n3930), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4958 (.d(n3931), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4959 (.d(n3932), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4960 (.d(n3933), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4961 (.d(n3934), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4962 (.d(n3935), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4963 (.d(n3936), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4964 (.d(n3937), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4965 (.d(n3938), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4966 (.d(n3939), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4967 (.d(n3940), .clk(clk), .s(1'b0), .r(rst), .q(\regs[9] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4968 (.d(n3941), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [31]));   // regs.v(41)
    VERIFIC_DFFRS i4969 (.d(n3942), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [30]));   // regs.v(41)
    VERIFIC_DFFRS i4970 (.d(n3943), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [29]));   // regs.v(41)
    VERIFIC_DFFRS i4971 (.d(n3944), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [28]));   // regs.v(41)
    VERIFIC_DFFRS i4972 (.d(n3945), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [27]));   // regs.v(41)
    VERIFIC_DFFRS i4973 (.d(n3946), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [26]));   // regs.v(41)
    VERIFIC_DFFRS i4974 (.d(n3947), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [25]));   // regs.v(41)
    VERIFIC_DFFRS i4975 (.d(n3948), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [24]));   // regs.v(41)
    VERIFIC_DFFRS i4976 (.d(n3949), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [23]));   // regs.v(41)
    VERIFIC_DFFRS i4977 (.d(n3950), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [22]));   // regs.v(41)
    VERIFIC_DFFRS i4978 (.d(n3951), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [21]));   // regs.v(41)
    VERIFIC_DFFRS i4979 (.d(n3952), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [20]));   // regs.v(41)
    VERIFIC_DFFRS i4980 (.d(n3953), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [19]));   // regs.v(41)
    VERIFIC_DFFRS i4981 (.d(n3954), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [18]));   // regs.v(41)
    VERIFIC_DFFRS i4982 (.d(n3955), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [17]));   // regs.v(41)
    VERIFIC_DFFRS i4983 (.d(n3956), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [16]));   // regs.v(41)
    VERIFIC_DFFRS i4984 (.d(n3957), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [15]));   // regs.v(41)
    VERIFIC_DFFRS i4985 (.d(n3958), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [14]));   // regs.v(41)
    VERIFIC_DFFRS i4986 (.d(n3959), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [13]));   // regs.v(41)
    VERIFIC_DFFRS i4987 (.d(n3960), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [12]));   // regs.v(41)
    VERIFIC_DFFRS i4988 (.d(n3961), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [11]));   // regs.v(41)
    VERIFIC_DFFRS i4989 (.d(n3962), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [10]));   // regs.v(41)
    VERIFIC_DFFRS i4990 (.d(n3963), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [9]));   // regs.v(41)
    VERIFIC_DFFRS i4991 (.d(n3964), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [8]));   // regs.v(41)
    VERIFIC_DFFRS i4992 (.d(n3965), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [7]));   // regs.v(41)
    VERIFIC_DFFRS i4993 (.d(n3966), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [6]));   // regs.v(41)
    VERIFIC_DFFRS i4994 (.d(n3967), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [5]));   // regs.v(41)
    VERIFIC_DFFRS i4995 (.d(n3968), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [4]));   // regs.v(41)
    VERIFIC_DFFRS i4996 (.d(n3969), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [3]));   // regs.v(41)
    VERIFIC_DFFRS i4997 (.d(n3970), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [2]));   // regs.v(41)
    VERIFIC_DFFRS i4998 (.d(n3971), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [1]));   // regs.v(41)
    VERIFIC_DFFRS i4999 (.d(n3972), .clk(clk), .s(1'b0), .r(rst), .q(\regs[8] [0]));   // regs.v(41)
    VERIFIC_DFFRS i5000 (.d(n3973), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [31]));   // regs.v(41)
    VERIFIC_DFFRS i5001 (.d(n3974), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [30]));   // regs.v(41)
    VERIFIC_DFFRS i5002 (.d(n3975), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [29]));   // regs.v(41)
    VERIFIC_DFFRS i5003 (.d(n3976), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [28]));   // regs.v(41)
    VERIFIC_DFFRS i5004 (.d(n3977), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [27]));   // regs.v(41)
    VERIFIC_DFFRS i5005 (.d(n3978), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [26]));   // regs.v(41)
    VERIFIC_DFFRS i5006 (.d(n3979), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [25]));   // regs.v(41)
    VERIFIC_DFFRS i5007 (.d(n3980), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [24]));   // regs.v(41)
    VERIFIC_DFFRS i5008 (.d(n3981), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [23]));   // regs.v(41)
    VERIFIC_DFFRS i5009 (.d(n3982), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [22]));   // regs.v(41)
    VERIFIC_DFFRS i5010 (.d(n3983), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [21]));   // regs.v(41)
    VERIFIC_DFFRS i5011 (.d(n3984), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [20]));   // regs.v(41)
    VERIFIC_DFFRS i5012 (.d(n3985), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [19]));   // regs.v(41)
    VERIFIC_DFFRS i5013 (.d(n3986), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [18]));   // regs.v(41)
    VERIFIC_DFFRS i5014 (.d(n3987), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [17]));   // regs.v(41)
    VERIFIC_DFFRS i5015 (.d(n3988), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [16]));   // regs.v(41)
    VERIFIC_DFFRS i5016 (.d(n3989), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [15]));   // regs.v(41)
    VERIFIC_DFFRS i5017 (.d(n3990), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [14]));   // regs.v(41)
    VERIFIC_DFFRS i5018 (.d(n3991), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [13]));   // regs.v(41)
    VERIFIC_DFFRS i5019 (.d(n3992), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [12]));   // regs.v(41)
    VERIFIC_DFFRS i5020 (.d(n3993), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [11]));   // regs.v(41)
    VERIFIC_DFFRS i5021 (.d(n3994), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [10]));   // regs.v(41)
    VERIFIC_DFFRS i5022 (.d(n3995), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [9]));   // regs.v(41)
    VERIFIC_DFFRS i5023 (.d(n3996), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [8]));   // regs.v(41)
    VERIFIC_DFFRS i5024 (.d(n3997), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [7]));   // regs.v(41)
    VERIFIC_DFFRS i5025 (.d(n3998), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [6]));   // regs.v(41)
    VERIFIC_DFFRS i5026 (.d(n3999), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [5]));   // regs.v(41)
    VERIFIC_DFFRS i5027 (.d(n4000), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [4]));   // regs.v(41)
    VERIFIC_DFFRS i5028 (.d(n4001), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [3]));   // regs.v(41)
    VERIFIC_DFFRS i5029 (.d(n4002), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [2]));   // regs.v(41)
    VERIFIC_DFFRS i5030 (.d(n4003), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [1]));   // regs.v(41)
    VERIFIC_DFFRS i5031 (.d(n4004), .clk(clk), .s(1'b0), .r(rst), .q(\regs[7] [0]));   // regs.v(41)
    VERIFIC_DFFRS i5032 (.d(n4005), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [31]));   // regs.v(41)
    VERIFIC_DFFRS i5033 (.d(n4006), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [30]));   // regs.v(41)
    VERIFIC_DFFRS i5034 (.d(n4007), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [29]));   // regs.v(41)
    VERIFIC_DFFRS i5035 (.d(n4008), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [28]));   // regs.v(41)
    VERIFIC_DFFRS i5036 (.d(n4009), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [27]));   // regs.v(41)
    VERIFIC_DFFRS i5037 (.d(n4010), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [26]));   // regs.v(41)
    VERIFIC_DFFRS i5038 (.d(n4011), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [25]));   // regs.v(41)
    VERIFIC_DFFRS i5039 (.d(n4012), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [24]));   // regs.v(41)
    VERIFIC_DFFRS i5040 (.d(n4013), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [23]));   // regs.v(41)
    VERIFIC_DFFRS i5041 (.d(n4014), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [22]));   // regs.v(41)
    VERIFIC_DFFRS i5042 (.d(n4015), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [21]));   // regs.v(41)
    VERIFIC_DFFRS i5043 (.d(n4016), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [20]));   // regs.v(41)
    VERIFIC_DFFRS i5044 (.d(n4017), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [19]));   // regs.v(41)
    VERIFIC_DFFRS i5045 (.d(n4018), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [18]));   // regs.v(41)
    VERIFIC_DFFRS i5046 (.d(n4019), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [17]));   // regs.v(41)
    VERIFIC_DFFRS i5047 (.d(n4020), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [16]));   // regs.v(41)
    VERIFIC_DFFRS i5048 (.d(n4021), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [15]));   // regs.v(41)
    VERIFIC_DFFRS i5049 (.d(n4022), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [14]));   // regs.v(41)
    VERIFIC_DFFRS i5050 (.d(n4023), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [13]));   // regs.v(41)
    VERIFIC_DFFRS i5051 (.d(n4024), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [12]));   // regs.v(41)
    VERIFIC_DFFRS i5052 (.d(n4025), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [11]));   // regs.v(41)
    VERIFIC_DFFRS i5053 (.d(n4026), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [10]));   // regs.v(41)
    VERIFIC_DFFRS i5054 (.d(n4027), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [9]));   // regs.v(41)
    VERIFIC_DFFRS i5055 (.d(n4028), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [8]));   // regs.v(41)
    VERIFIC_DFFRS i5056 (.d(n4029), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [7]));   // regs.v(41)
    VERIFIC_DFFRS i5057 (.d(n4030), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [6]));   // regs.v(41)
    VERIFIC_DFFRS i5058 (.d(n4031), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [5]));   // regs.v(41)
    VERIFIC_DFFRS i5059 (.d(n4032), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [4]));   // regs.v(41)
    VERIFIC_DFFRS i5060 (.d(n4033), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [3]));   // regs.v(41)
    VERIFIC_DFFRS i5061 (.d(n4034), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [2]));   // regs.v(41)
    VERIFIC_DFFRS i5062 (.d(n4035), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [1]));   // regs.v(41)
    VERIFIC_DFFRS i5063 (.d(n4036), .clk(clk), .s(1'b0), .r(rst), .q(\regs[6] [0]));   // regs.v(41)
    VERIFIC_DFFRS i5064 (.d(n4037), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [31]));   // regs.v(41)
    VERIFIC_DFFRS i5065 (.d(n4038), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [30]));   // regs.v(41)
    VERIFIC_DFFRS i5066 (.d(n4039), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [29]));   // regs.v(41)
    VERIFIC_DFFRS i5067 (.d(n4040), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [28]));   // regs.v(41)
    VERIFIC_DFFRS i5068 (.d(n4041), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [27]));   // regs.v(41)
    VERIFIC_DFFRS i5069 (.d(n4042), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [26]));   // regs.v(41)
    VERIFIC_DFFRS i5070 (.d(n4043), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [25]));   // regs.v(41)
    VERIFIC_DFFRS i5071 (.d(n4044), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [24]));   // regs.v(41)
    VERIFIC_DFFRS i5072 (.d(n4045), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [23]));   // regs.v(41)
    VERIFIC_DFFRS i5073 (.d(n4046), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [22]));   // regs.v(41)
    VERIFIC_DFFRS i5074 (.d(n4047), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [21]));   // regs.v(41)
    VERIFIC_DFFRS i5075 (.d(n4048), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [20]));   // regs.v(41)
    VERIFIC_DFFRS i5076 (.d(n4049), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [19]));   // regs.v(41)
    VERIFIC_DFFRS i5077 (.d(n4050), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [18]));   // regs.v(41)
    VERIFIC_DFFRS i5078 (.d(n4051), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [17]));   // regs.v(41)
    VERIFIC_DFFRS i5079 (.d(n4052), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [16]));   // regs.v(41)
    VERIFIC_DFFRS i5080 (.d(n4053), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [15]));   // regs.v(41)
    VERIFIC_DFFRS i5081 (.d(n4054), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [14]));   // regs.v(41)
    VERIFIC_DFFRS i5082 (.d(n4055), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [13]));   // regs.v(41)
    VERIFIC_DFFRS i5083 (.d(n4056), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [12]));   // regs.v(41)
    VERIFIC_DFFRS i5084 (.d(n4057), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [11]));   // regs.v(41)
    VERIFIC_DFFRS i5085 (.d(n4058), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [10]));   // regs.v(41)
    VERIFIC_DFFRS i5086 (.d(n4059), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [9]));   // regs.v(41)
    VERIFIC_DFFRS i5087 (.d(n4060), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [8]));   // regs.v(41)
    VERIFIC_DFFRS i5088 (.d(n4061), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [7]));   // regs.v(41)
    VERIFIC_DFFRS i5089 (.d(n4062), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [6]));   // regs.v(41)
    VERIFIC_DFFRS i5090 (.d(n4063), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [5]));   // regs.v(41)
    VERIFIC_DFFRS i5091 (.d(n4064), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [4]));   // regs.v(41)
    VERIFIC_DFFRS i5092 (.d(n4065), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [3]));   // regs.v(41)
    VERIFIC_DFFRS i5093 (.d(n4066), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [2]));   // regs.v(41)
    VERIFIC_DFFRS i5094 (.d(n4067), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [1]));   // regs.v(41)
    VERIFIC_DFFRS i5095 (.d(n4068), .clk(clk), .s(1'b0), .r(rst), .q(\regs[5] [0]));   // regs.v(41)
    VERIFIC_DFFRS i5096 (.d(n4069), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [31]));   // regs.v(41)
    VERIFIC_DFFRS i5097 (.d(n4070), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [30]));   // regs.v(41)
    VERIFIC_DFFRS i5098 (.d(n4071), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [29]));   // regs.v(41)
    VERIFIC_DFFRS i5099 (.d(n4072), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [28]));   // regs.v(41)
    VERIFIC_DFFRS i5100 (.d(n4073), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [27]));   // regs.v(41)
    VERIFIC_DFFRS i5101 (.d(n4074), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [26]));   // regs.v(41)
    VERIFIC_DFFRS i5102 (.d(n4075), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [25]));   // regs.v(41)
    VERIFIC_DFFRS i5103 (.d(n4076), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [24]));   // regs.v(41)
    VERIFIC_DFFRS i5104 (.d(n4077), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [23]));   // regs.v(41)
    VERIFIC_DFFRS i5105 (.d(n4078), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [22]));   // regs.v(41)
    VERIFIC_DFFRS i5106 (.d(n4079), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [21]));   // regs.v(41)
    VERIFIC_DFFRS i5107 (.d(n4080), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [20]));   // regs.v(41)
    VERIFIC_DFFRS i5108 (.d(n4081), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [19]));   // regs.v(41)
    VERIFIC_DFFRS i5109 (.d(n4082), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [18]));   // regs.v(41)
    VERIFIC_DFFRS i5110 (.d(n4083), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [17]));   // regs.v(41)
    VERIFIC_DFFRS i5111 (.d(n4084), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [16]));   // regs.v(41)
    VERIFIC_DFFRS i5112 (.d(n4085), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [15]));   // regs.v(41)
    VERIFIC_DFFRS i5113 (.d(n4086), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [14]));   // regs.v(41)
    VERIFIC_DFFRS i5114 (.d(n4087), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [13]));   // regs.v(41)
    VERIFIC_DFFRS i5115 (.d(n4088), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [12]));   // regs.v(41)
    VERIFIC_DFFRS i5116 (.d(n4089), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [11]));   // regs.v(41)
    VERIFIC_DFFRS i5117 (.d(n4090), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [10]));   // regs.v(41)
    VERIFIC_DFFRS i5118 (.d(n4091), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [9]));   // regs.v(41)
    VERIFIC_DFFRS i5119 (.d(n4092), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [8]));   // regs.v(41)
    VERIFIC_DFFRS i5120 (.d(n4093), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [7]));   // regs.v(41)
    VERIFIC_DFFRS i5121 (.d(n4094), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [6]));   // regs.v(41)
    VERIFIC_DFFRS i5122 (.d(n4095), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [5]));   // regs.v(41)
    VERIFIC_DFFRS i5123 (.d(n4096), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [4]));   // regs.v(41)
    VERIFIC_DFFRS i5124 (.d(n4097), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [3]));   // regs.v(41)
    VERIFIC_DFFRS i5125 (.d(n4098), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [2]));   // regs.v(41)
    VERIFIC_DFFRS i5126 (.d(n4099), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [1]));   // regs.v(41)
    VERIFIC_DFFRS i5127 (.d(n4100), .clk(clk), .s(1'b0), .r(rst), .q(\regs[4] [0]));   // regs.v(41)
    VERIFIC_DFFRS i5128 (.d(n4101), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [31]));   // regs.v(41)
    VERIFIC_DFFRS i5129 (.d(n4102), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [30]));   // regs.v(41)
    VERIFIC_DFFRS i5130 (.d(n4103), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [29]));   // regs.v(41)
    VERIFIC_DFFRS i5131 (.d(n4104), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [28]));   // regs.v(41)
    VERIFIC_DFFRS i5132 (.d(n4105), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [27]));   // regs.v(41)
    VERIFIC_DFFRS i5133 (.d(n4106), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [26]));   // regs.v(41)
    VERIFIC_DFFRS i5134 (.d(n4107), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [25]));   // regs.v(41)
    VERIFIC_DFFRS i5135 (.d(n4108), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [24]));   // regs.v(41)
    VERIFIC_DFFRS i5136 (.d(n4109), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [23]));   // regs.v(41)
    VERIFIC_DFFRS i5137 (.d(n4110), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [22]));   // regs.v(41)
    VERIFIC_DFFRS i5138 (.d(n4111), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [21]));   // regs.v(41)
    VERIFIC_DFFRS i5139 (.d(n4112), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [20]));   // regs.v(41)
    VERIFIC_DFFRS i5140 (.d(n4113), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [19]));   // regs.v(41)
    VERIFIC_DFFRS i5141 (.d(n4114), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [18]));   // regs.v(41)
    VERIFIC_DFFRS i5142 (.d(n4115), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [17]));   // regs.v(41)
    VERIFIC_DFFRS i5143 (.d(n4116), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [16]));   // regs.v(41)
    VERIFIC_DFFRS i5144 (.d(n4117), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [15]));   // regs.v(41)
    VERIFIC_DFFRS i5145 (.d(n4118), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [14]));   // regs.v(41)
    VERIFIC_DFFRS i5146 (.d(n4119), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [13]));   // regs.v(41)
    VERIFIC_DFFRS i5147 (.d(n4120), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [12]));   // regs.v(41)
    VERIFIC_DFFRS i5148 (.d(n4121), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [11]));   // regs.v(41)
    VERIFIC_DFFRS i5149 (.d(n4122), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [10]));   // regs.v(41)
    VERIFIC_DFFRS i5150 (.d(n4123), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [9]));   // regs.v(41)
    VERIFIC_DFFRS i5151 (.d(n4124), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [8]));   // regs.v(41)
    VERIFIC_DFFRS i5152 (.d(n4125), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [7]));   // regs.v(41)
    VERIFIC_DFFRS i5153 (.d(n4126), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [6]));   // regs.v(41)
    VERIFIC_DFFRS i5154 (.d(n4127), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [5]));   // regs.v(41)
    VERIFIC_DFFRS i5155 (.d(n4128), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [4]));   // regs.v(41)
    VERIFIC_DFFRS i5156 (.d(n4129), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [3]));   // regs.v(41)
    VERIFIC_DFFRS i5157 (.d(n4130), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [2]));   // regs.v(41)
    VERIFIC_DFFRS i5158 (.d(n4131), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [1]));   // regs.v(41)
    VERIFIC_DFFRS i5159 (.d(n4132), .clk(clk), .s(1'b0), .r(rst), .q(\regs[3] [0]));   // regs.v(41)
    VERIFIC_DFFRS i5160 (.d(n4133), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [31]));   // regs.v(41)
    VERIFIC_DFFRS i5161 (.d(n4134), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [30]));   // regs.v(41)
    VERIFIC_DFFRS i5162 (.d(n4135), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [29]));   // regs.v(41)
    VERIFIC_DFFRS i5163 (.d(n4136), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [28]));   // regs.v(41)
    VERIFIC_DFFRS i5164 (.d(n4137), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [27]));   // regs.v(41)
    VERIFIC_DFFRS i5165 (.d(n4138), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [26]));   // regs.v(41)
    VERIFIC_DFFRS i5166 (.d(n4139), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [25]));   // regs.v(41)
    VERIFIC_DFFRS i5167 (.d(n4140), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [24]));   // regs.v(41)
    VERIFIC_DFFRS i5168 (.d(n4141), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [23]));   // regs.v(41)
    VERIFIC_DFFRS i5169 (.d(n4142), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [22]));   // regs.v(41)
    VERIFIC_DFFRS i5170 (.d(n4143), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [21]));   // regs.v(41)
    VERIFIC_DFFRS i5171 (.d(n4144), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [20]));   // regs.v(41)
    VERIFIC_DFFRS i5172 (.d(n4145), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [19]));   // regs.v(41)
    VERIFIC_DFFRS i5173 (.d(n4146), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [18]));   // regs.v(41)
    VERIFIC_DFFRS i5174 (.d(n4147), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [17]));   // regs.v(41)
    VERIFIC_DFFRS i5175 (.d(n4148), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [16]));   // regs.v(41)
    VERIFIC_DFFRS i5176 (.d(n4149), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [15]));   // regs.v(41)
    VERIFIC_DFFRS i5177 (.d(n4150), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [14]));   // regs.v(41)
    VERIFIC_DFFRS i5178 (.d(n4151), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [13]));   // regs.v(41)
    VERIFIC_DFFRS i5179 (.d(n4152), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [12]));   // regs.v(41)
    VERIFIC_DFFRS i5180 (.d(n4153), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [11]));   // regs.v(41)
    VERIFIC_DFFRS i5181 (.d(n4154), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [10]));   // regs.v(41)
    VERIFIC_DFFRS i5182 (.d(n4155), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [9]));   // regs.v(41)
    VERIFIC_DFFRS i5183 (.d(n4156), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [8]));   // regs.v(41)
    VERIFIC_DFFRS i5184 (.d(n4157), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [7]));   // regs.v(41)
    VERIFIC_DFFRS i5185 (.d(n4158), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [6]));   // regs.v(41)
    VERIFIC_DFFRS i5186 (.d(n4159), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [5]));   // regs.v(41)
    VERIFIC_DFFRS i5187 (.d(n4160), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [4]));   // regs.v(41)
    VERIFIC_DFFRS i5188 (.d(n4161), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [3]));   // regs.v(41)
    VERIFIC_DFFRS i5189 (.d(n4162), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [2]));   // regs.v(41)
    VERIFIC_DFFRS i5190 (.d(n4163), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [1]));   // regs.v(41)
    VERIFIC_DFFRS i5191 (.d(n4164), .clk(clk), .s(1'b0), .r(rst), .q(\regs[2] [0]));   // regs.v(41)
    VERIFIC_DFFRS i5192 (.d(n4165), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [31]));   // regs.v(41)
    VERIFIC_DFFRS i5193 (.d(n4166), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [30]));   // regs.v(41)
    VERIFIC_DFFRS i5194 (.d(n4167), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [29]));   // regs.v(41)
    VERIFIC_DFFRS i5195 (.d(n4168), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [28]));   // regs.v(41)
    VERIFIC_DFFRS i5196 (.d(n4169), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [27]));   // regs.v(41)
    VERIFIC_DFFRS i5197 (.d(n4170), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [26]));   // regs.v(41)
    VERIFIC_DFFRS i5198 (.d(n4171), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [25]));   // regs.v(41)
    VERIFIC_DFFRS i5199 (.d(n4172), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [24]));   // regs.v(41)
    VERIFIC_DFFRS i5200 (.d(n4173), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [23]));   // regs.v(41)
    VERIFIC_DFFRS i5201 (.d(n4174), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [22]));   // regs.v(41)
    VERIFIC_DFFRS i5202 (.d(n4175), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [21]));   // regs.v(41)
    VERIFIC_DFFRS i5203 (.d(n4176), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [20]));   // regs.v(41)
    VERIFIC_DFFRS i5204 (.d(n4177), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [19]));   // regs.v(41)
    VERIFIC_DFFRS i5205 (.d(n4178), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [18]));   // regs.v(41)
    VERIFIC_DFFRS i5206 (.d(n4179), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [17]));   // regs.v(41)
    VERIFIC_DFFRS i5207 (.d(n4180), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [16]));   // regs.v(41)
    VERIFIC_DFFRS i5208 (.d(n4181), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [15]));   // regs.v(41)
    VERIFIC_DFFRS i5209 (.d(n4182), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [14]));   // regs.v(41)
    VERIFIC_DFFRS i5210 (.d(n4183), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [13]));   // regs.v(41)
    VERIFIC_DFFRS i5211 (.d(n4184), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [12]));   // regs.v(41)
    VERIFIC_DFFRS i5212 (.d(n4185), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [11]));   // regs.v(41)
    VERIFIC_DFFRS i5213 (.d(n4186), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [10]));   // regs.v(41)
    VERIFIC_DFFRS i5214 (.d(n4187), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [9]));   // regs.v(41)
    VERIFIC_DFFRS i5215 (.d(n4188), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [8]));   // regs.v(41)
    VERIFIC_DFFRS i5216 (.d(n4189), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [7]));   // regs.v(41)
    VERIFIC_DFFRS i5217 (.d(n4190), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [6]));   // regs.v(41)
    VERIFIC_DFFRS i5218 (.d(n4191), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [5]));   // regs.v(41)
    VERIFIC_DFFRS i5219 (.d(n4192), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [4]));   // regs.v(41)
    VERIFIC_DFFRS i5220 (.d(n4193), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [3]));   // regs.v(41)
    VERIFIC_DFFRS i5221 (.d(n4194), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [2]));   // regs.v(41)
    VERIFIC_DFFRS i5222 (.d(n4195), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [1]));   // regs.v(41)
    VERIFIC_DFFRS i5223 (.d(n4196), .clk(clk), .s(1'b0), .r(rst), .q(\regs[1] [0]));   // regs.v(41)
    VERIFIC_DFFRS i5224 (.d(n4197), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [31]));   // regs.v(41)
    VERIFIC_DFFRS i5225 (.d(n4198), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [30]));   // regs.v(41)
    VERIFIC_DFFRS i5226 (.d(n4199), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [29]));   // regs.v(41)
    VERIFIC_DFFRS i5227 (.d(n4200), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [28]));   // regs.v(41)
    VERIFIC_DFFRS i5228 (.d(n4201), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [27]));   // regs.v(41)
    VERIFIC_DFFRS i5229 (.d(n4202), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [26]));   // regs.v(41)
    VERIFIC_DFFRS i5230 (.d(n4203), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [25]));   // regs.v(41)
    VERIFIC_DFFRS i5231 (.d(n4204), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [24]));   // regs.v(41)
    VERIFIC_DFFRS i5232 (.d(n4205), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [23]));   // regs.v(41)
    VERIFIC_DFFRS i5233 (.d(n4206), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [22]));   // regs.v(41)
    VERIFIC_DFFRS i5234 (.d(n4207), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [21]));   // regs.v(41)
    VERIFIC_DFFRS i5235 (.d(n4208), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [20]));   // regs.v(41)
    VERIFIC_DFFRS i5236 (.d(n4209), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [19]));   // regs.v(41)
    VERIFIC_DFFRS i5237 (.d(n4210), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [18]));   // regs.v(41)
    VERIFIC_DFFRS i5238 (.d(n4211), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [17]));   // regs.v(41)
    VERIFIC_DFFRS i5239 (.d(n4212), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [16]));   // regs.v(41)
    VERIFIC_DFFRS i5240 (.d(n4213), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [15]));   // regs.v(41)
    VERIFIC_DFFRS i5241 (.d(n4214), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [14]));   // regs.v(41)
    VERIFIC_DFFRS i5242 (.d(n4215), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [13]));   // regs.v(41)
    VERIFIC_DFFRS i5243 (.d(n4216), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [12]));   // regs.v(41)
    VERIFIC_DFFRS i5244 (.d(n4217), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [11]));   // regs.v(41)
    VERIFIC_DFFRS i5245 (.d(n4218), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [10]));   // regs.v(41)
    VERIFIC_DFFRS i5246 (.d(n4219), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [9]));   // regs.v(41)
    VERIFIC_DFFRS i5247 (.d(n4220), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [8]));   // regs.v(41)
    VERIFIC_DFFRS i5248 (.d(n4221), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [7]));   // regs.v(41)
    VERIFIC_DFFRS i5249 (.d(n4222), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [6]));   // regs.v(41)
    VERIFIC_DFFRS i5250 (.d(n4223), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [5]));   // regs.v(41)
    VERIFIC_DFFRS i5251 (.d(n4224), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [4]));   // regs.v(41)
    VERIFIC_DFFRS i5252 (.d(n4225), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [3]));   // regs.v(41)
    VERIFIC_DFFRS i5253 (.d(n4226), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [2]));   // regs.v(41)
    VERIFIC_DFFRS i5254 (.d(n4227), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [1]));   // regs.v(41)
    VERIFIC_DFFRS i5255 (.d(n4228), .clk(clk), .s(1'b0), .r(rst), .q(\regs[0] [0]));   // regs.v(41)
    VERIFIC_DFFRS i4232 (.d(n4294), .clk(clk), .s(1'b0), .r(rst), .q(pcout[31]));   // regs.v(41)
    
endmodule

//
// Verific Verilog Description of OPERATOR Mux_5u_32u
//

module Mux_5u_32u (sel, data, o);
    input [4:0]sel;
    input [31:0]data;
    output o;
    assign o = data[sel];
    
endmodule

//
// Verific Verilog Description of OPERATOR Decoder_5
//

module Decoder_5 (i, o);
    input [4:0]i;
    output [31:0]o;
    reg [31:0]o;
    always @(i) begin
    o = 0;
    o[i] = 1'b1;
    end
    
endmodule

//
// Verific Verilog Description of OPERATOR add_32u_32u
//

module add_32u_32u (cin, a, b, o, cout);
    input cin;
    input [31:0]a;
    input [31:0]b;
    output [31:0]o;
    output cout;
    assign {cout, o} = a + b + cin;
    
endmodule

//
// Verific Verilog Description of PRIMITIVE VERIFIC_DFFRS
//

module VERIFIC_DFFRS (d, clk, s, r, q);
    input d;
    input clk;
    input s;
    input r;
    output q;
    reg q ;
    always @(posedge clk or posedge s or posedge r) begin
        if (s) q = 1'b1;
        else if (r) q = 1'b0;
        else q = d;
    end
    
endmodule

//
// Verific Verilog Description of module insn_decoder
//

module insn_decoder (e_a, e_b, e_alu_op, e_is_cond, e_cond, e_write_flags, 
            e_swp, m_a1, m_a2, m_r1_op, m_r2_op, r_a1, r_a2, r_op, 
            d_pass, d_pcincr, r_r1_addr, r_r2_addr, r_read, word, 
            r1, r2, hazard, rst, clk);   // insn_decoder.v(89)
    output [31:0]e_a;   // insn_decoder.v(90)
    output [31:0]e_b;   // insn_decoder.v(90)
    output [7:0]e_alu_op;   // insn_decoder.v(91)
    output e_is_cond;   // insn_decoder.v(95)
    output [3:0]e_cond;   // insn_decoder.v(92)
    output [3:0]e_write_flags;   // insn_decoder.v(93)
    output e_swp;   // insn_decoder.v(94)
    output [31:0]m_a1;   // insn_decoder.v(97)
    output [31:0]m_a2;   // insn_decoder.v(97)
    output [3:0]m_r1_op;   // insn_decoder.v(98)
    output [3:0]m_r2_op;   // insn_decoder.v(98)
    output [4:0]r_a1;   // insn_decoder.v(100)
    output [4:0]r_a2;   // insn_decoder.v(100)
    output [3:0]r_op;   // insn_decoder.v(101)
    output d_pass;   // insn_decoder.v(103)
    output d_pcincr;   // insn_decoder.v(104)
    output [4:0]r_r1_addr;   // insn_decoder.v(106)
    output [4:0]r_r2_addr;   // insn_decoder.v(106)
    output [1:0]r_read;   // insn_decoder.v(107)
    input [31:0]word;   // insn_decoder.v(109)
    input [31:0]r1;   // insn_decoder.v(110)
    input [31:0]r2;   // insn_decoder.v(110)
    input hazard;   // insn_decoder.v(111)
    input rst;   // insn_decoder.v(112)
    input clk;   // insn_decoder.v(112)
    
    wire [7:0]state1;   // insn_decoder.v(114)
    wire fetch;   // insn_decoder.v(115)
    wire reg_fetch;   // insn_decoder.v(116)
    wire [3:0]delay_counter;   // insn_decoder.v(117)
    wire [2:0]imm_action;   // insn_decoder.v(118)
    wire [7:0]old_state1_imm;   // insn_decoder.v(120)
    wire old_pass_imm;   // insn_decoder.v(121)
    wire old_fetch_imm;   // insn_decoder.v(121)
    wire old_pcincr_imm;   // insn_decoder.v(121)
    wire [1:0]r_to_mem;   // insn_decoder.v(122)
    wire [7:0]old_state1_hz;   // insn_decoder.v(123)
    wire old_pass_hz;   // insn_decoder.v(124)
    wire old_fetch_hz;   // insn_decoder.v(124)
    wire old_pcincr_hz;   // insn_decoder.v(124)
    wire set_delay;   // insn_decoder.v(125)
    wire [3:0]cond;   // insn_decoder.v(128)
    wire [4:0]reg_a_addr;   // insn_decoder.v(130)
    wire [4:0]reg_b_addr;   // insn_decoder.v(130)
    wire [4:0]reg_c_addr;   // insn_decoder.v(131)
    wire [4:0]reg_d_addr;   // insn_decoder.v(131)
    
    wire n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
        n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, 
        n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
        n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, 
        n52, n53, n57, n59, n60, n65, n68, n69, n70, n71, 
        n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
        n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, 
        n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, 
        n102, n103, n104, n105, n106, n107, n108, n109, n110, 
        n111, n112, n113, n114, n115, n116, n117, n118, n119, 
        n120, n121, n122, n123, n124, n125, n126, n127, n128, 
        n129, n130, n131, n132, n133, n134, n135, n136, n137, 
        n138, n139, n140, n141, n142, n143, n144, n145, n146, 
        n147, n148, n149, n150, n151, n152, n153, n154, n155, 
        n156, n157, n158, n159, n160, n161, n162, n163, n164, 
        n165, n166, n167, n168, n169, n170, n171, n172, n173, 
        n174, n175, n176, n177, n178, n179, n180, n181, n182, 
        n183, n184, n185, n186, n187, n188, n189, n190, n191, 
        n192, n193, n194, n195, n196, n197, n198, n199, n200, 
        n201, n202, n203, n204, n205, n206, n207, n208, n209, 
        n210, n211, n212, n213, n214, n215, n216, n217, n218, 
        n219, n220, n221, n222, n223, n224, n225, n226, n227, 
        n228, n229, n230, n231, n232, n233, n234, n235, n236, 
        n237, n238, n239, n240, n241, n242, n243, n244, n245, 
        n246, n247, n248, n249, n250, n251, n252, n253, n254, 
        n255, n256, n257, n258, n259, n260, n261, n262, n263, 
        n264, n265, n266, n267, n268, n269, n270, n271, n272, 
        n273, n274, n275, n276, n277, n278, n279, n280, n281, 
        n282, n283, n284, n285, n286, n287, n288, n289, n290, 
        n291, n292, n293, n294, n295, n296, n297, n298, n299, 
        n300, n301, n302, n303, n304, n305, n306, n307, n308, 
        n309, n310, n311, n312, n313, n314, n315, n316, n317, 
        n318, n319, n320, n321, n322, n323, n324, n325, n326, 
        n327, n328, n329, n330, n331, n332, n333, n334, n335, 
        n336, n337, n338, n339, n340, n341, n342, n343, n344, 
        n345, n346, n347, n348, n349, n350, n351, n352, n353, 
        n354, n355, n356, n357, n358, n359, n360, n361, n362, 
        n363, n364, n365, n366, n367, n368, n369, n370, n371, 
        n372, n373, n374, n375, n376, n377, n378, n379, n380, 
        n381, n382, n383, n384, n385, n386, n387, n388, n391, 
        n395, n396, n397, n398, n399, n400, n401, n402, n403, 
        n404, n405, n406, n407, n408, n409, n410, n411, n412, 
        n413, n414, n415, n416, n417, n418, n419, n420, n421, 
        n422, n423, n424, n425, n426, n427, n428, n429, n430, 
        n431, n432, n433, n434, n435, n436, n437, n438, n439, 
        n440, n441, n442, n443, n444, n445, n446, n447, n448, 
        n449, n450, n451, n452, n453, n454, n455, n456, n457, 
        n458, n459, n460, n461, n462, n463, n464, n465, n466, 
        n467, n468, n469, n470, n471, n472, n473, n474, n475, 
        n476, n477, n478, n479, n480, n481, n482, n483, n484, 
        n485, n486, n487, n488, n489, n490, n491, n492, n494, 
        n495, n496, n497, n498, n499, n500, n501, n502, n503, 
        n504, n505, n506, n507, n508, n509, n510, n511, n512, 
        n513, n514, n515, n516, n517, n518, n519, n520, n521, 
        n522, n523, n524, n525, n526, n527, n528, n531, n532, 
        n533, n536, n539, n546, n547, n548, n551, n554, n558, 
        n561, n565, n569, n574, n575, n576, n579, n582, n586, 
        n589, n593, n597, n602, n605, n609, n613, n618, n622, 
        n627, n632, n638, n639, n640, n643, n644, n651, n655, 
        n656, n657, n658, n659, n660, n661, n662, n663, n664, 
        n665, n666, n667, n668, n669, n670, n671, n672, n673, 
        n674, n675, n676, n677, n678, n679, n680, n681, n682, 
        n683, n684, n685, n686, n687, n688, n689, n690, n691, 
        n692, n693, n694, n695, n696, n697, n698, n699, n700, 
        n701, n702, n703, n704, n705, n706, n707, n708, n709, 
        n710, n711, n712, n713, n714, n715, n716, n717, n718, 
        n719, n720, n721, n722, n723, n724, n725, n726, n727, 
        n728, n729, n730, n731, n732, n733, n734, n735, n736, 
        n737, n738, n739, n740, n741, n742, n743, n744, n745, 
        n746, n747, n748, n749, n750, n751, n752, n753, n754, 
        n755, n756, n757, n758, n759, n760, n761, n762, n763, 
        n764, n765, n766, n767, n768, n769, n770, n771, n772, 
        n774, n776, n777, n778, n780, n781, n782, n784, n785, 
        n786, n788, n789, n790, n792, n793, n794, n796, n797, 
        n799, n802, n805, n808, n809, n810, n812, n816, n820, 
        n824, n827, n828, n830, n832, n833, n835, n836, n837, 
        n839, n840, n842, n843, n845, n848, n851, n853, n854, 
        n855, n857, n858, n859, n861, n862, n863, n865, n866, 
        n867, n869, n872, n874, n875, n876, n878, n879, n880, 
        n881, n882, n886, n890, n894, n898, n899, n900, n901, 
        n902, n906, n910, n913, n917, n918, n919, n920, n923, 
        n926, n929, n932, n933, n934, n936, n939, n941, n942, 
        n943, n944, n945, n948, n951, n954, n957, n958, n959, 
        n960, n963, n966, n969, n972, n975, n978, n981, n984, 
        n987, n990, n993, n996, n999, n1002, n1005, n1008, n1011, 
        n1014, n1017, n1020, n1023, n1026, n1029, n1032, n1035, 
        n1038, n1041, n1044, n1047, n1050, n1053, n1054, n1056, 
        n1057, n1059, n1062, n1064, n1065, n1068, n1071, n1074, 
        n1077, n1080, n1083, n1084, n1086, n1089, n1092, n1095, 
        n1097, n1099, n1101, n1103, n1105, n1107, n1109, n1111, 
        n1113, n1115, n1117, n1119, n1121, n1123, n1125, n1127, 
        n1129, n1131, n1133, n1135, n1137, n1139, n1141, n1143, 
        n1145, n1147, n1149, n1151, n1153, n1155, n1157, n1159, 
        n1161, n1163, n1165, n1167, n1169, n1171, n1173, n1175, 
        n1177, n1179, n1181, n1183, n1185, n1187, n1189, n1191, 
        n1193, n1195, n1197, n1199, n1201, n1203, n1205, n1207, 
        n1209, n1211, n1213, n1215, n1217, n1219, n1221, n1223, 
        n1224, n1225, n1227, n1229, n1231, n1233, n1235, n1237, 
        n1239, n1241, n1243, n1245, n1247, n1249, n1251, n1253, 
        n1255, n1257, n1259, n1261, n1263, n1265, n1267, n1269, 
        n1271, n1273, n1275, n1277, n1279, n1281, n1283, n1285, 
        n1287, n1288, n1289, n1291, n1292, n1293, n1294, n1295, 
        n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1304, 
        n1305, n1306, n1308, n1311, n1312, n1313, n1314, n1316, 
        n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, 
        n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, 
        n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, 
        n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, 
        n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
        n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, 
        n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, 
        n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, 
        n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, 
        n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
        n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, 
        n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, 
        n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, 
        n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, 
        n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
        n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, 
        n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, 
        n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, 
        n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, 
        n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, 
        n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, 
        n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, 
        n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, 
        n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, 
        n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
        n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, 
        n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, 
        n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, 
        n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, 
        n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
        n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, 
        n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, 
        n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, 
        n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, 
        n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, 
        n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, 
        n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, 
        n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, 
        n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, 
        n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, 
        n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, 
        n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, 
        n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, 
        n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, 
        n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
        n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, 
        n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, 
        n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, 
        n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, 
        n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
        n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, 
        n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, 
        n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, 
        n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, 
        n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, 
        n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, 
        n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, 
        n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, 
        n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, 
        n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, 
        n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, 
        n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, 
        n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
        n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, 
        n2073, n2074, n2075, n2076, n2082, n2083, n2084, n2085, 
        n2086, n2092, n2093, n2094, n2095, n2096, n2102, n2103, 
        n2104, n2105, n2106, n2112, n2113, n2114, n2115, n2116;
    
    assign n12 = fetch ? word[24] : cond[3];   // insn_decoder.v(185)
    assign n13 = fetch ? word[23] : cond[2];   // insn_decoder.v(185)
    assign n14 = fetch ? word[22] : cond[1];   // insn_decoder.v(185)
    assign n15 = fetch ? word[21] : cond[0];   // insn_decoder.v(185)
    assign n16 = fetch ? word[20] : reg_a_addr[4];   // insn_decoder.v(185)
    assign n17 = fetch ? word[19] : reg_a_addr[3];   // insn_decoder.v(185)
    assign n18 = fetch ? word[18] : reg_a_addr[2];   // insn_decoder.v(185)
    assign n19 = fetch ? word[17] : reg_a_addr[1];   // insn_decoder.v(185)
    assign n20 = fetch ? word[16] : reg_a_addr[0];   // insn_decoder.v(185)
    assign n21 = fetch ? word[15] : reg_b_addr[4];   // insn_decoder.v(185)
    assign n22 = fetch ? word[14] : reg_b_addr[3];   // insn_decoder.v(185)
    assign n23 = fetch ? word[13] : reg_b_addr[2];   // insn_decoder.v(185)
    assign n24 = fetch ? word[12] : reg_b_addr[1];   // insn_decoder.v(185)
    assign n25 = fetch ? word[11] : reg_b_addr[0];   // insn_decoder.v(185)
    assign n26 = fetch ? word[10] : reg_c_addr[4];   // insn_decoder.v(185)
    assign n27 = fetch ? word[9] : reg_c_addr[3];   // insn_decoder.v(185)
    assign n28 = fetch ? word[8] : reg_c_addr[2];   // insn_decoder.v(185)
    assign n29 = fetch ? word[7] : reg_c_addr[1];   // insn_decoder.v(185)
    assign n30 = fetch ? word[6] : reg_c_addr[0];   // insn_decoder.v(185)
    assign n31 = fetch ? word[5] : reg_d_addr[4];   // insn_decoder.v(185)
    assign n32 = fetch ? word[4] : reg_d_addr[3];   // insn_decoder.v(185)
    assign n33 = fetch ? word[3] : reg_d_addr[2];   // insn_decoder.v(185)
    assign n34 = fetch ? word[2] : reg_d_addr[1];   // insn_decoder.v(185)
    assign n35 = fetch ? word[1] : reg_d_addr[0];   // insn_decoder.v(185)
    assign n36 = fetch ? 1'b0 : imm_action[2];   // insn_decoder.v(185)
    assign n37 = fetch ? word[5] : imm_action[1];   // insn_decoder.v(185)
    assign n38 = fetch ? word[4] : imm_action[0];   // insn_decoder.v(185)
    assign n39 = fetch ? 1'b0 : state1[7];   // insn_decoder.v(185)
    assign n40 = fetch ? word[31] : state1[6];   // insn_decoder.v(185)
    assign n41 = fetch ? word[30] : state1[5];   // insn_decoder.v(185)
    assign n42 = fetch ? word[29] : state1[4];   // insn_decoder.v(185)
    assign n43 = fetch ? word[28] : state1[3];   // insn_decoder.v(185)
    assign n44 = fetch ? word[27] : state1[2];   // insn_decoder.v(185)
    assign n45 = fetch ? word[26] : state1[1];   // insn_decoder.v(185)
    assign n46 = fetch ? word[25] : state1[0];   // insn_decoder.v(185)
    assign n47 = fetch ? 1'b1 : d_pcincr;   // insn_decoder.v(185)
    assign n48 = fetch ? 1'b1 : d_pass;   // insn_decoder.v(185)
    assign n49 = fetch ? 1'b1 : reg_fetch;   // insn_decoder.v(185)
    not (n50, imm_action[0]) ;   // insn_decoder.v(520)
    nor (n51, imm_action[2], imm_action[1], n50) ;   // insn_decoder.v(520)
    not (n52, imm_action[1]) ;   // insn_decoder.v(521)
    nor (n53, imm_action[2], n52, imm_action[0]) ;   // insn_decoder.v(521)
    nor (n391, imm_action[2], n52, n50) ;   // insn_decoder.v(521)
    or (n57, n53, n391) ;   // insn_decoder.v(521)
    not (n59, imm_action[2]) ;   // insn_decoder.v(522)
    nor (n60, n59, n52, imm_action[0]) ;   // insn_decoder.v(522)
    nor (n395, n59, n52, n50) ;   // insn_decoder.v(522)
    or (n65, n60, n395) ;   // insn_decoder.v(522)
    nor (n68, n59, imm_action[1], n50) ;   // insn_decoder.v(523)
    assign n69 = n68 ? word[31] : m_a2[31];   // insn_decoder.v(523)
    assign n70 = n68 ? word[30] : m_a2[30];   // insn_decoder.v(523)
    assign n71 = n68 ? word[29] : m_a2[29];   // insn_decoder.v(523)
    assign n72 = n68 ? word[28] : m_a2[28];   // insn_decoder.v(523)
    assign n73 = n68 ? word[27] : m_a2[27];   // insn_decoder.v(523)
    assign n74 = n68 ? word[26] : m_a2[26];   // insn_decoder.v(523)
    assign n75 = n68 ? word[25] : m_a2[25];   // insn_decoder.v(523)
    assign n76 = n68 ? word[24] : m_a2[24];   // insn_decoder.v(523)
    assign n77 = n68 ? word[23] : m_a2[23];   // insn_decoder.v(523)
    assign n78 = n68 ? word[22] : m_a2[22];   // insn_decoder.v(523)
    assign n79 = n68 ? word[21] : m_a2[21];   // insn_decoder.v(523)
    assign n80 = n68 ? word[20] : m_a2[20];   // insn_decoder.v(523)
    assign n81 = n68 ? word[19] : m_a2[19];   // insn_decoder.v(523)
    assign n82 = n68 ? word[18] : m_a2[18];   // insn_decoder.v(523)
    assign n83 = n68 ? word[17] : m_a2[17];   // insn_decoder.v(523)
    assign n84 = n68 ? word[16] : m_a2[16];   // insn_decoder.v(523)
    assign n85 = n68 ? word[15] : m_a2[15];   // insn_decoder.v(523)
    assign n86 = n68 ? word[14] : m_a2[14];   // insn_decoder.v(523)
    assign n87 = n68 ? word[13] : m_a2[13];   // insn_decoder.v(523)
    assign n88 = n68 ? word[12] : m_a2[12];   // insn_decoder.v(523)
    assign n89 = n68 ? word[11] : m_a2[11];   // insn_decoder.v(523)
    assign n90 = n68 ? word[10] : m_a2[10];   // insn_decoder.v(523)
    assign n91 = n68 ? word[9] : m_a2[9];   // insn_decoder.v(523)
    assign n92 = n68 ? word[8] : m_a2[8];   // insn_decoder.v(523)
    assign n93 = n68 ? word[7] : m_a2[7];   // insn_decoder.v(523)
    assign n94 = n68 ? word[6] : m_a2[6];   // insn_decoder.v(523)
    assign n95 = n68 ? word[5] : m_a2[5];   // insn_decoder.v(523)
    assign n96 = n68 ? word[4] : m_a2[4];   // insn_decoder.v(523)
    assign n97 = n68 ? word[3] : m_a2[3];   // insn_decoder.v(523)
    assign n98 = n68 ? word[2] : m_a2[2];   // insn_decoder.v(523)
    assign n99 = n68 ? word[1] : m_a2[1];   // insn_decoder.v(523)
    assign n100 = n68 ? word[0] : m_a2[0];   // insn_decoder.v(523)
    assign n101 = n65 ? word[31] : m_a1[31];   // insn_decoder.v(523)
    assign n102 = n65 ? word[30] : m_a1[30];   // insn_decoder.v(523)
    assign n103 = n65 ? word[29] : m_a1[29];   // insn_decoder.v(523)
    assign n104 = n65 ? word[28] : m_a1[28];   // insn_decoder.v(523)
    assign n105 = n65 ? word[27] : m_a1[27];   // insn_decoder.v(523)
    assign n106 = n65 ? word[26] : m_a1[26];   // insn_decoder.v(523)
    assign n107 = n65 ? word[25] : m_a1[25];   // insn_decoder.v(523)
    assign n108 = n65 ? word[24] : m_a1[24];   // insn_decoder.v(523)
    assign n109 = n65 ? word[23] : m_a1[23];   // insn_decoder.v(523)
    assign n110 = n65 ? word[22] : m_a1[22];   // insn_decoder.v(523)
    assign n111 = n65 ? word[21] : m_a1[21];   // insn_decoder.v(523)
    assign n112 = n65 ? word[20] : m_a1[20];   // insn_decoder.v(523)
    assign n113 = n65 ? word[19] : m_a1[19];   // insn_decoder.v(523)
    assign n114 = n65 ? word[18] : m_a1[18];   // insn_decoder.v(523)
    assign n115 = n65 ? word[17] : m_a1[17];   // insn_decoder.v(523)
    assign n116 = n65 ? word[16] : m_a1[16];   // insn_decoder.v(523)
    assign n117 = n65 ? word[15] : m_a1[15];   // insn_decoder.v(523)
    assign n118 = n65 ? word[14] : m_a1[14];   // insn_decoder.v(523)
    assign n119 = n65 ? word[13] : m_a1[13];   // insn_decoder.v(523)
    assign n120 = n65 ? word[12] : m_a1[12];   // insn_decoder.v(523)
    assign n121 = n65 ? word[11] : m_a1[11];   // insn_decoder.v(523)
    assign n122 = n65 ? word[10] : m_a1[10];   // insn_decoder.v(523)
    assign n123 = n65 ? word[9] : m_a1[9];   // insn_decoder.v(523)
    assign n124 = n65 ? word[8] : m_a1[8];   // insn_decoder.v(523)
    assign n125 = n65 ? word[7] : m_a1[7];   // insn_decoder.v(523)
    assign n126 = n65 ? word[6] : m_a1[6];   // insn_decoder.v(523)
    assign n127 = n65 ? word[5] : m_a1[5];   // insn_decoder.v(523)
    assign n128 = n65 ? word[4] : m_a1[4];   // insn_decoder.v(523)
    assign n129 = n65 ? word[3] : m_a1[3];   // insn_decoder.v(523)
    assign n130 = n65 ? word[2] : m_a1[2];   // insn_decoder.v(523)
    assign n131 = n65 ? word[1] : m_a1[1];   // insn_decoder.v(523)
    assign n132 = n65 ? word[0] : m_a1[0];   // insn_decoder.v(523)
    assign n133 = n65 ? m_a2[31] : n69;   // insn_decoder.v(523)
    assign n134 = n65 ? m_a2[30] : n70;   // insn_decoder.v(523)
    assign n135 = n65 ? m_a2[29] : n71;   // insn_decoder.v(523)
    assign n136 = n65 ? m_a2[28] : n72;   // insn_decoder.v(523)
    assign n137 = n65 ? m_a2[27] : n73;   // insn_decoder.v(523)
    assign n138 = n65 ? m_a2[26] : n74;   // insn_decoder.v(523)
    assign n139 = n65 ? m_a2[25] : n75;   // insn_decoder.v(523)
    assign n140 = n65 ? m_a2[24] : n76;   // insn_decoder.v(523)
    assign n141 = n65 ? m_a2[23] : n77;   // insn_decoder.v(523)
    assign n142 = n65 ? m_a2[22] : n78;   // insn_decoder.v(523)
    assign n143 = n65 ? m_a2[21] : n79;   // insn_decoder.v(523)
    assign n144 = n65 ? m_a2[20] : n80;   // insn_decoder.v(523)
    assign n145 = n65 ? m_a2[19] : n81;   // insn_decoder.v(523)
    assign n146 = n65 ? m_a2[18] : n82;   // insn_decoder.v(523)
    assign n147 = n65 ? m_a2[17] : n83;   // insn_decoder.v(523)
    assign n148 = n65 ? m_a2[16] : n84;   // insn_decoder.v(523)
    assign n149 = n65 ? m_a2[15] : n85;   // insn_decoder.v(523)
    assign n150 = n65 ? m_a2[14] : n86;   // insn_decoder.v(523)
    assign n151 = n65 ? m_a2[13] : n87;   // insn_decoder.v(523)
    assign n152 = n65 ? m_a2[12] : n88;   // insn_decoder.v(523)
    assign n153 = n65 ? m_a2[11] : n89;   // insn_decoder.v(523)
    assign n154 = n65 ? m_a2[10] : n90;   // insn_decoder.v(523)
    assign n155 = n65 ? m_a2[9] : n91;   // insn_decoder.v(523)
    assign n156 = n65 ? m_a2[8] : n92;   // insn_decoder.v(523)
    assign n157 = n65 ? m_a2[7] : n93;   // insn_decoder.v(523)
    assign n158 = n65 ? m_a2[6] : n94;   // insn_decoder.v(523)
    assign n159 = n65 ? m_a2[5] : n95;   // insn_decoder.v(523)
    assign n160 = n65 ? m_a2[4] : n96;   // insn_decoder.v(523)
    assign n161 = n65 ? m_a2[3] : n97;   // insn_decoder.v(523)
    assign n162 = n65 ? m_a2[2] : n98;   // insn_decoder.v(523)
    assign n163 = n65 ? m_a2[1] : n99;   // insn_decoder.v(523)
    assign n164 = n65 ? m_a2[0] : n100;   // insn_decoder.v(523)
    assign n165 = n57 ? word[31] : e_a[31];   // insn_decoder.v(522)
    assign n166 = n57 ? word[30] : e_a[30];   // insn_decoder.v(522)
    assign n167 = n57 ? word[29] : e_a[29];   // insn_decoder.v(522)
    assign n168 = n57 ? word[28] : e_a[28];   // insn_decoder.v(522)
    assign n169 = n57 ? word[27] : e_a[27];   // insn_decoder.v(522)
    assign n170 = n57 ? word[26] : e_a[26];   // insn_decoder.v(522)
    assign n171 = n57 ? word[25] : e_a[25];   // insn_decoder.v(522)
    assign n172 = n57 ? word[24] : e_a[24];   // insn_decoder.v(522)
    assign n173 = n57 ? word[23] : e_a[23];   // insn_decoder.v(522)
    assign n174 = n57 ? word[22] : e_a[22];   // insn_decoder.v(522)
    assign n175 = n57 ? word[21] : e_a[21];   // insn_decoder.v(522)
    assign n176 = n57 ? word[20] : e_a[20];   // insn_decoder.v(522)
    assign n177 = n57 ? word[19] : e_a[19];   // insn_decoder.v(522)
    assign n178 = n57 ? word[18] : e_a[18];   // insn_decoder.v(522)
    assign n179 = n57 ? word[17] : e_a[17];   // insn_decoder.v(522)
    assign n180 = n57 ? word[16] : e_a[16];   // insn_decoder.v(522)
    assign n181 = n57 ? word[15] : e_a[15];   // insn_decoder.v(522)
    assign n182 = n57 ? word[14] : e_a[14];   // insn_decoder.v(522)
    assign n183 = n57 ? word[13] : e_a[13];   // insn_decoder.v(522)
    assign n184 = n57 ? word[12] : e_a[12];   // insn_decoder.v(522)
    assign n185 = n57 ? word[11] : e_a[11];   // insn_decoder.v(522)
    assign n186 = n57 ? word[10] : e_a[10];   // insn_decoder.v(522)
    assign n187 = n57 ? word[9] : e_a[9];   // insn_decoder.v(522)
    assign n188 = n57 ? word[8] : e_a[8];   // insn_decoder.v(522)
    assign n189 = n57 ? word[7] : e_a[7];   // insn_decoder.v(522)
    assign n190 = n57 ? word[6] : e_a[6];   // insn_decoder.v(522)
    assign n191 = n57 ? word[5] : e_a[5];   // insn_decoder.v(522)
    assign n192 = n57 ? word[4] : e_a[4];   // insn_decoder.v(522)
    assign n193 = n57 ? word[3] : e_a[3];   // insn_decoder.v(522)
    assign n194 = n57 ? word[2] : e_a[2];   // insn_decoder.v(522)
    assign n195 = n57 ? word[1] : e_a[1];   // insn_decoder.v(522)
    assign n196 = n57 ? word[0] : e_a[0];   // insn_decoder.v(522)
    assign n197 = n57 ? m_a1[31] : n101;   // insn_decoder.v(522)
    assign n198 = n57 ? m_a1[30] : n102;   // insn_decoder.v(522)
    assign n199 = n57 ? m_a1[29] : n103;   // insn_decoder.v(522)
    assign n200 = n57 ? m_a1[28] : n104;   // insn_decoder.v(522)
    assign n201 = n57 ? m_a1[27] : n105;   // insn_decoder.v(522)
    assign n202 = n57 ? m_a1[26] : n106;   // insn_decoder.v(522)
    assign n203 = n57 ? m_a1[25] : n107;   // insn_decoder.v(522)
    assign n204 = n57 ? m_a1[24] : n108;   // insn_decoder.v(522)
    assign n205 = n57 ? m_a1[23] : n109;   // insn_decoder.v(522)
    assign n206 = n57 ? m_a1[22] : n110;   // insn_decoder.v(522)
    assign n207 = n57 ? m_a1[21] : n111;   // insn_decoder.v(522)
    assign n208 = n57 ? m_a1[20] : n112;   // insn_decoder.v(522)
    assign n209 = n57 ? m_a1[19] : n113;   // insn_decoder.v(522)
    assign n210 = n57 ? m_a1[18] : n114;   // insn_decoder.v(522)
    assign n211 = n57 ? m_a1[17] : n115;   // insn_decoder.v(522)
    assign n212 = n57 ? m_a1[16] : n116;   // insn_decoder.v(522)
    assign n213 = n57 ? m_a1[15] : n117;   // insn_decoder.v(522)
    assign n214 = n57 ? m_a1[14] : n118;   // insn_decoder.v(522)
    assign n215 = n57 ? m_a1[13] : n119;   // insn_decoder.v(522)
    assign n216 = n57 ? m_a1[12] : n120;   // insn_decoder.v(522)
    assign n217 = n57 ? m_a1[11] : n121;   // insn_decoder.v(522)
    assign n218 = n57 ? m_a1[10] : n122;   // insn_decoder.v(522)
    assign n219 = n57 ? m_a1[9] : n123;   // insn_decoder.v(522)
    assign n220 = n57 ? m_a1[8] : n124;   // insn_decoder.v(522)
    assign n221 = n57 ? m_a1[7] : n125;   // insn_decoder.v(522)
    assign n222 = n57 ? m_a1[6] : n126;   // insn_decoder.v(522)
    assign n223 = n57 ? m_a1[5] : n127;   // insn_decoder.v(522)
    assign n224 = n57 ? m_a1[4] : n128;   // insn_decoder.v(522)
    assign n225 = n57 ? m_a1[3] : n129;   // insn_decoder.v(522)
    assign n226 = n57 ? m_a1[2] : n130;   // insn_decoder.v(522)
    assign n227 = n57 ? m_a1[1] : n131;   // insn_decoder.v(522)
    assign n228 = n57 ? m_a1[0] : n132;   // insn_decoder.v(522)
    assign n229 = n57 ? m_a2[31] : n133;   // insn_decoder.v(522)
    assign n230 = n57 ? m_a2[30] : n134;   // insn_decoder.v(522)
    assign n231 = n57 ? m_a2[29] : n135;   // insn_decoder.v(522)
    assign n232 = n57 ? m_a2[28] : n136;   // insn_decoder.v(522)
    assign n233 = n57 ? m_a2[27] : n137;   // insn_decoder.v(522)
    assign n234 = n57 ? m_a2[26] : n138;   // insn_decoder.v(522)
    assign n235 = n57 ? m_a2[25] : n139;   // insn_decoder.v(522)
    assign n236 = n57 ? m_a2[24] : n140;   // insn_decoder.v(522)
    assign n237 = n57 ? m_a2[23] : n141;   // insn_decoder.v(522)
    assign n238 = n57 ? m_a2[22] : n142;   // insn_decoder.v(522)
    assign n239 = n57 ? m_a2[21] : n143;   // insn_decoder.v(522)
    assign n240 = n57 ? m_a2[20] : n144;   // insn_decoder.v(522)
    assign n241 = n57 ? m_a2[19] : n145;   // insn_decoder.v(522)
    assign n242 = n57 ? m_a2[18] : n146;   // insn_decoder.v(522)
    assign n243 = n57 ? m_a2[17] : n147;   // insn_decoder.v(522)
    assign n244 = n57 ? m_a2[16] : n148;   // insn_decoder.v(522)
    assign n245 = n57 ? m_a2[15] : n149;   // insn_decoder.v(522)
    assign n246 = n57 ? m_a2[14] : n150;   // insn_decoder.v(522)
    assign n247 = n57 ? m_a2[13] : n151;   // insn_decoder.v(522)
    assign n248 = n57 ? m_a2[12] : n152;   // insn_decoder.v(522)
    assign n249 = n57 ? m_a2[11] : n153;   // insn_decoder.v(522)
    assign n250 = n57 ? m_a2[10] : n154;   // insn_decoder.v(522)
    assign n251 = n57 ? m_a2[9] : n155;   // insn_decoder.v(522)
    assign n252 = n57 ? m_a2[8] : n156;   // insn_decoder.v(522)
    assign n253 = n57 ? m_a2[7] : n157;   // insn_decoder.v(522)
    assign n254 = n57 ? m_a2[6] : n158;   // insn_decoder.v(522)
    assign n255 = n57 ? m_a2[5] : n159;   // insn_decoder.v(522)
    assign n256 = n57 ? m_a2[4] : n160;   // insn_decoder.v(522)
    assign n257 = n57 ? m_a2[3] : n161;   // insn_decoder.v(522)
    assign n258 = n57 ? m_a2[2] : n162;   // insn_decoder.v(522)
    assign n259 = n57 ? m_a2[1] : n163;   // insn_decoder.v(522)
    assign n260 = n57 ? m_a2[0] : n164;   // insn_decoder.v(522)
    assign n261 = n51 ? word[31] : e_b[31];   // insn_decoder.v(521)
    assign n262 = n51 ? word[30] : e_b[30];   // insn_decoder.v(521)
    assign n263 = n51 ? word[29] : e_b[29];   // insn_decoder.v(521)
    assign n264 = n51 ? word[28] : e_b[28];   // insn_decoder.v(521)
    assign n265 = n51 ? word[27] : e_b[27];   // insn_decoder.v(521)
    assign n266 = n51 ? word[26] : e_b[26];   // insn_decoder.v(521)
    assign n267 = n51 ? word[25] : e_b[25];   // insn_decoder.v(521)
    assign n268 = n51 ? word[24] : e_b[24];   // insn_decoder.v(521)
    assign n269 = n51 ? word[23] : e_b[23];   // insn_decoder.v(521)
    assign n270 = n51 ? word[22] : e_b[22];   // insn_decoder.v(521)
    assign n271 = n51 ? word[21] : e_b[21];   // insn_decoder.v(521)
    assign n272 = n51 ? word[20] : e_b[20];   // insn_decoder.v(521)
    assign n273 = n51 ? word[19] : e_b[19];   // insn_decoder.v(521)
    assign n274 = n51 ? word[18] : e_b[18];   // insn_decoder.v(521)
    assign n275 = n51 ? word[17] : e_b[17];   // insn_decoder.v(521)
    assign n276 = n51 ? word[16] : e_b[16];   // insn_decoder.v(521)
    assign n277 = n51 ? word[15] : e_b[15];   // insn_decoder.v(521)
    assign n278 = n51 ? word[14] : e_b[14];   // insn_decoder.v(521)
    assign n279 = n51 ? word[13] : e_b[13];   // insn_decoder.v(521)
    assign n280 = n51 ? word[12] : e_b[12];   // insn_decoder.v(521)
    assign n281 = n51 ? word[11] : e_b[11];   // insn_decoder.v(521)
    assign n282 = n51 ? word[10] : e_b[10];   // insn_decoder.v(521)
    assign n283 = n51 ? word[9] : e_b[9];   // insn_decoder.v(521)
    assign n284 = n51 ? word[8] : e_b[8];   // insn_decoder.v(521)
    assign n285 = n51 ? word[7] : e_b[7];   // insn_decoder.v(521)
    assign n286 = n51 ? word[6] : e_b[6];   // insn_decoder.v(521)
    assign n287 = n51 ? word[5] : e_b[5];   // insn_decoder.v(521)
    assign n288 = n51 ? word[4] : e_b[4];   // insn_decoder.v(521)
    assign n289 = n51 ? word[3] : e_b[3];   // insn_decoder.v(521)
    assign n290 = n51 ? word[2] : e_b[2];   // insn_decoder.v(521)
    assign n291 = n51 ? word[1] : e_b[1];   // insn_decoder.v(521)
    assign n292 = n51 ? word[0] : e_b[0];   // insn_decoder.v(521)
    assign n293 = n51 ? e_a[31] : n165;   // insn_decoder.v(521)
    assign n294 = n51 ? e_a[30] : n166;   // insn_decoder.v(521)
    assign n295 = n51 ? e_a[29] : n167;   // insn_decoder.v(521)
    assign n296 = n51 ? e_a[28] : n168;   // insn_decoder.v(521)
    assign n297 = n51 ? e_a[27] : n169;   // insn_decoder.v(521)
    assign n298 = n51 ? e_a[26] : n170;   // insn_decoder.v(521)
    assign n299 = n51 ? e_a[25] : n171;   // insn_decoder.v(521)
    assign n300 = n51 ? e_a[24] : n172;   // insn_decoder.v(521)
    assign n301 = n51 ? e_a[23] : n173;   // insn_decoder.v(521)
    assign n302 = n51 ? e_a[22] : n174;   // insn_decoder.v(521)
    assign n303 = n51 ? e_a[21] : n175;   // insn_decoder.v(521)
    assign n304 = n51 ? e_a[20] : n176;   // insn_decoder.v(521)
    assign n305 = n51 ? e_a[19] : n177;   // insn_decoder.v(521)
    assign n306 = n51 ? e_a[18] : n178;   // insn_decoder.v(521)
    assign n307 = n51 ? e_a[17] : n179;   // insn_decoder.v(521)
    assign n308 = n51 ? e_a[16] : n180;   // insn_decoder.v(521)
    assign n309 = n51 ? e_a[15] : n181;   // insn_decoder.v(521)
    assign n310 = n51 ? e_a[14] : n182;   // insn_decoder.v(521)
    assign n311 = n51 ? e_a[13] : n183;   // insn_decoder.v(521)
    assign n312 = n51 ? e_a[12] : n184;   // insn_decoder.v(521)
    assign n313 = n51 ? e_a[11] : n185;   // insn_decoder.v(521)
    assign n314 = n51 ? e_a[10] : n186;   // insn_decoder.v(521)
    assign n315 = n51 ? e_a[9] : n187;   // insn_decoder.v(521)
    assign n316 = n51 ? e_a[8] : n188;   // insn_decoder.v(521)
    assign n317 = n51 ? e_a[7] : n189;   // insn_decoder.v(521)
    assign n318 = n51 ? e_a[6] : n190;   // insn_decoder.v(521)
    assign n319 = n51 ? e_a[5] : n191;   // insn_decoder.v(521)
    assign n320 = n51 ? e_a[4] : n192;   // insn_decoder.v(521)
    assign n321 = n51 ? e_a[3] : n193;   // insn_decoder.v(521)
    assign n322 = n51 ? e_a[2] : n194;   // insn_decoder.v(521)
    assign n323 = n51 ? e_a[1] : n195;   // insn_decoder.v(521)
    assign n324 = n51 ? e_a[0] : n196;   // insn_decoder.v(521)
    assign n325 = n51 ? m_a1[31] : n197;   // insn_decoder.v(521)
    assign n326 = n51 ? m_a1[30] : n198;   // insn_decoder.v(521)
    assign n327 = n51 ? m_a1[29] : n199;   // insn_decoder.v(521)
    assign n328 = n51 ? m_a1[28] : n200;   // insn_decoder.v(521)
    assign n329 = n51 ? m_a1[27] : n201;   // insn_decoder.v(521)
    assign n330 = n51 ? m_a1[26] : n202;   // insn_decoder.v(521)
    assign n331 = n51 ? m_a1[25] : n203;   // insn_decoder.v(521)
    assign n332 = n51 ? m_a1[24] : n204;   // insn_decoder.v(521)
    assign n333 = n51 ? m_a1[23] : n205;   // insn_decoder.v(521)
    assign n334 = n51 ? m_a1[22] : n206;   // insn_decoder.v(521)
    assign n335 = n51 ? m_a1[21] : n207;   // insn_decoder.v(521)
    assign n336 = n51 ? m_a1[20] : n208;   // insn_decoder.v(521)
    assign n337 = n51 ? m_a1[19] : n209;   // insn_decoder.v(521)
    assign n338 = n51 ? m_a1[18] : n210;   // insn_decoder.v(521)
    assign n339 = n51 ? m_a1[17] : n211;   // insn_decoder.v(521)
    assign n340 = n51 ? m_a1[16] : n212;   // insn_decoder.v(521)
    assign n341 = n51 ? m_a1[15] : n213;   // insn_decoder.v(521)
    assign n342 = n51 ? m_a1[14] : n214;   // insn_decoder.v(521)
    assign n343 = n51 ? m_a1[13] : n215;   // insn_decoder.v(521)
    assign n344 = n51 ? m_a1[12] : n216;   // insn_decoder.v(521)
    assign n345 = n51 ? m_a1[11] : n217;   // insn_decoder.v(521)
    assign n346 = n51 ? m_a1[10] : n218;   // insn_decoder.v(521)
    assign n347 = n51 ? m_a1[9] : n219;   // insn_decoder.v(521)
    assign n348 = n51 ? m_a1[8] : n220;   // insn_decoder.v(521)
    assign n349 = n51 ? m_a1[7] : n221;   // insn_decoder.v(521)
    assign n350 = n51 ? m_a1[6] : n222;   // insn_decoder.v(521)
    assign n351 = n51 ? m_a1[5] : n223;   // insn_decoder.v(521)
    assign n352 = n51 ? m_a1[4] : n224;   // insn_decoder.v(521)
    assign n353 = n51 ? m_a1[3] : n225;   // insn_decoder.v(521)
    assign n354 = n51 ? m_a1[2] : n226;   // insn_decoder.v(521)
    assign n355 = n51 ? m_a1[1] : n227;   // insn_decoder.v(521)
    assign n356 = n51 ? m_a1[0] : n228;   // insn_decoder.v(521)
    assign n357 = n51 ? m_a2[31] : n229;   // insn_decoder.v(521)
    assign n358 = n51 ? m_a2[30] : n230;   // insn_decoder.v(521)
    assign n359 = n51 ? m_a2[29] : n231;   // insn_decoder.v(521)
    assign n360 = n51 ? m_a2[28] : n232;   // insn_decoder.v(521)
    assign n361 = n51 ? m_a2[27] : n233;   // insn_decoder.v(521)
    assign n362 = n51 ? m_a2[26] : n234;   // insn_decoder.v(521)
    assign n363 = n51 ? m_a2[25] : n235;   // insn_decoder.v(521)
    assign n364 = n51 ? m_a2[24] : n236;   // insn_decoder.v(521)
    assign n365 = n51 ? m_a2[23] : n237;   // insn_decoder.v(521)
    assign n366 = n51 ? m_a2[22] : n238;   // insn_decoder.v(521)
    assign n367 = n51 ? m_a2[21] : n239;   // insn_decoder.v(521)
    assign n368 = n51 ? m_a2[20] : n240;   // insn_decoder.v(521)
    assign n369 = n51 ? m_a2[19] : n241;   // insn_decoder.v(521)
    assign n370 = n51 ? m_a2[18] : n242;   // insn_decoder.v(521)
    assign n371 = n51 ? m_a2[17] : n243;   // insn_decoder.v(521)
    assign n372 = n51 ? m_a2[16] : n244;   // insn_decoder.v(521)
    assign n373 = n51 ? m_a2[15] : n245;   // insn_decoder.v(521)
    assign n374 = n51 ? m_a2[14] : n246;   // insn_decoder.v(521)
    assign n375 = n51 ? m_a2[13] : n247;   // insn_decoder.v(521)
    assign n376 = n51 ? m_a2[12] : n248;   // insn_decoder.v(521)
    assign n377 = n51 ? m_a2[11] : n249;   // insn_decoder.v(521)
    assign n378 = n51 ? m_a2[10] : n250;   // insn_decoder.v(521)
    assign n379 = n51 ? m_a2[9] : n251;   // insn_decoder.v(521)
    assign n380 = n51 ? m_a2[8] : n252;   // insn_decoder.v(521)
    assign n381 = n51 ? m_a2[7] : n253;   // insn_decoder.v(521)
    assign n382 = n51 ? m_a2[6] : n254;   // insn_decoder.v(521)
    assign n383 = n51 ? m_a2[5] : n255;   // insn_decoder.v(521)
    assign n384 = n51 ? m_a2[4] : n256;   // insn_decoder.v(521)
    assign n385 = n51 ? m_a2[3] : n257;   // insn_decoder.v(521)
    assign n386 = n51 ? m_a2[2] : n258;   // insn_decoder.v(521)
    assign n387 = n51 ? m_a2[1] : n259;   // insn_decoder.v(521)
    assign n388 = n51 ? m_a2[0] : n260;   // insn_decoder.v(521)
    assign n396 = n395 ? word[31] : m_a2[31];   // insn_decoder.v(527)
    assign n397 = n395 ? word[30] : m_a2[30];   // insn_decoder.v(527)
    assign n398 = n395 ? word[29] : m_a2[29];   // insn_decoder.v(527)
    assign n399 = n395 ? word[28] : m_a2[28];   // insn_decoder.v(527)
    assign n400 = n395 ? word[27] : m_a2[27];   // insn_decoder.v(527)
    assign n401 = n395 ? word[26] : m_a2[26];   // insn_decoder.v(527)
    assign n402 = n395 ? word[25] : m_a2[25];   // insn_decoder.v(527)
    assign n403 = n395 ? word[24] : m_a2[24];   // insn_decoder.v(527)
    assign n404 = n395 ? word[23] : m_a2[23];   // insn_decoder.v(527)
    assign n405 = n395 ? word[22] : m_a2[22];   // insn_decoder.v(527)
    assign n406 = n395 ? word[21] : m_a2[21];   // insn_decoder.v(527)
    assign n407 = n395 ? word[20] : m_a2[20];   // insn_decoder.v(527)
    assign n408 = n395 ? word[19] : m_a2[19];   // insn_decoder.v(527)
    assign n409 = n395 ? word[18] : m_a2[18];   // insn_decoder.v(527)
    assign n410 = n395 ? word[17] : m_a2[17];   // insn_decoder.v(527)
    assign n411 = n395 ? word[16] : m_a2[16];   // insn_decoder.v(527)
    assign n412 = n395 ? word[15] : m_a2[15];   // insn_decoder.v(527)
    assign n413 = n395 ? word[14] : m_a2[14];   // insn_decoder.v(527)
    assign n414 = n395 ? word[13] : m_a2[13];   // insn_decoder.v(527)
    assign n415 = n395 ? word[12] : m_a2[12];   // insn_decoder.v(527)
    assign n416 = n395 ? word[11] : m_a2[11];   // insn_decoder.v(527)
    assign n417 = n395 ? word[10] : m_a2[10];   // insn_decoder.v(527)
    assign n418 = n395 ? word[9] : m_a2[9];   // insn_decoder.v(527)
    assign n419 = n395 ? word[8] : m_a2[8];   // insn_decoder.v(527)
    assign n420 = n395 ? word[7] : m_a2[7];   // insn_decoder.v(527)
    assign n421 = n395 ? word[6] : m_a2[6];   // insn_decoder.v(527)
    assign n422 = n395 ? word[5] : m_a2[5];   // insn_decoder.v(527)
    assign n423 = n395 ? word[4] : m_a2[4];   // insn_decoder.v(527)
    assign n424 = n395 ? word[3] : m_a2[3];   // insn_decoder.v(527)
    assign n425 = n395 ? word[2] : m_a2[2];   // insn_decoder.v(527)
    assign n426 = n395 ? word[1] : m_a2[1];   // insn_decoder.v(527)
    assign n427 = n395 ? word[0] : m_a2[0];   // insn_decoder.v(527)
    assign n428 = n391 ? word[31] : e_b[31];   // insn_decoder.v(527)
    assign n429 = n391 ? word[30] : e_b[30];   // insn_decoder.v(527)
    assign n430 = n391 ? word[29] : e_b[29];   // insn_decoder.v(527)
    assign n431 = n391 ? word[28] : e_b[28];   // insn_decoder.v(527)
    assign n432 = n391 ? word[27] : e_b[27];   // insn_decoder.v(527)
    assign n433 = n391 ? word[26] : e_b[26];   // insn_decoder.v(527)
    assign n434 = n391 ? word[25] : e_b[25];   // insn_decoder.v(527)
    assign n435 = n391 ? word[24] : e_b[24];   // insn_decoder.v(527)
    assign n436 = n391 ? word[23] : e_b[23];   // insn_decoder.v(527)
    assign n437 = n391 ? word[22] : e_b[22];   // insn_decoder.v(527)
    assign n438 = n391 ? word[21] : e_b[21];   // insn_decoder.v(527)
    assign n439 = n391 ? word[20] : e_b[20];   // insn_decoder.v(527)
    assign n440 = n391 ? word[19] : e_b[19];   // insn_decoder.v(527)
    assign n441 = n391 ? word[18] : e_b[18];   // insn_decoder.v(527)
    assign n442 = n391 ? word[17] : e_b[17];   // insn_decoder.v(527)
    assign n443 = n391 ? word[16] : e_b[16];   // insn_decoder.v(527)
    assign n444 = n391 ? word[15] : e_b[15];   // insn_decoder.v(527)
    assign n445 = n391 ? word[14] : e_b[14];   // insn_decoder.v(527)
    assign n446 = n391 ? word[13] : e_b[13];   // insn_decoder.v(527)
    assign n447 = n391 ? word[12] : e_b[12];   // insn_decoder.v(527)
    assign n448 = n391 ? word[11] : e_b[11];   // insn_decoder.v(527)
    assign n449 = n391 ? word[10] : e_b[10];   // insn_decoder.v(527)
    assign n450 = n391 ? word[9] : e_b[9];   // insn_decoder.v(527)
    assign n451 = n391 ? word[8] : e_b[8];   // insn_decoder.v(527)
    assign n452 = n391 ? word[7] : e_b[7];   // insn_decoder.v(527)
    assign n453 = n391 ? word[6] : e_b[6];   // insn_decoder.v(527)
    assign n454 = n391 ? word[5] : e_b[5];   // insn_decoder.v(527)
    assign n455 = n391 ? word[4] : e_b[4];   // insn_decoder.v(527)
    assign n456 = n391 ? word[3] : e_b[3];   // insn_decoder.v(527)
    assign n457 = n391 ? word[2] : e_b[2];   // insn_decoder.v(527)
    assign n458 = n391 ? word[1] : e_b[1];   // insn_decoder.v(527)
    assign n459 = n391 ? word[0] : e_b[0];   // insn_decoder.v(527)
    assign n460 = n391 ? m_a2[31] : n396;   // insn_decoder.v(527)
    assign n461 = n391 ? m_a2[30] : n397;   // insn_decoder.v(527)
    assign n462 = n391 ? m_a2[29] : n398;   // insn_decoder.v(527)
    assign n463 = n391 ? m_a2[28] : n399;   // insn_decoder.v(527)
    assign n464 = n391 ? m_a2[27] : n400;   // insn_decoder.v(527)
    assign n465 = n391 ? m_a2[26] : n401;   // insn_decoder.v(527)
    assign n466 = n391 ? m_a2[25] : n402;   // insn_decoder.v(527)
    assign n467 = n391 ? m_a2[24] : n403;   // insn_decoder.v(527)
    assign n468 = n391 ? m_a2[23] : n404;   // insn_decoder.v(527)
    assign n469 = n391 ? m_a2[22] : n405;   // insn_decoder.v(527)
    assign n470 = n391 ? m_a2[21] : n406;   // insn_decoder.v(527)
    assign n471 = n391 ? m_a2[20] : n407;   // insn_decoder.v(527)
    assign n472 = n391 ? m_a2[19] : n408;   // insn_decoder.v(527)
    assign n473 = n391 ? m_a2[18] : n409;   // insn_decoder.v(527)
    assign n474 = n391 ? m_a2[17] : n410;   // insn_decoder.v(527)
    assign n475 = n391 ? m_a2[16] : n411;   // insn_decoder.v(527)
    assign n476 = n391 ? m_a2[15] : n412;   // insn_decoder.v(527)
    assign n477 = n391 ? m_a2[14] : n413;   // insn_decoder.v(527)
    assign n478 = n391 ? m_a2[13] : n414;   // insn_decoder.v(527)
    assign n479 = n391 ? m_a2[12] : n415;   // insn_decoder.v(527)
    assign n480 = n391 ? m_a2[11] : n416;   // insn_decoder.v(527)
    assign n481 = n391 ? m_a2[10] : n417;   // insn_decoder.v(527)
    assign n482 = n391 ? m_a2[9] : n418;   // insn_decoder.v(527)
    assign n483 = n391 ? m_a2[8] : n419;   // insn_decoder.v(527)
    assign n484 = n391 ? m_a2[7] : n420;   // insn_decoder.v(527)
    assign n485 = n391 ? m_a2[6] : n421;   // insn_decoder.v(527)
    assign n486 = n391 ? m_a2[5] : n422;   // insn_decoder.v(527)
    assign n487 = n391 ? m_a2[4] : n423;   // insn_decoder.v(527)
    assign n488 = n391 ? m_a2[3] : n424;   // insn_decoder.v(527)
    assign n489 = n391 ? m_a2[2] : n425;   // insn_decoder.v(527)
    assign n490 = n391 ? m_a2[1] : n426;   // insn_decoder.v(527)
    assign n491 = n391 ? m_a2[0] : n427;   // insn_decoder.v(527)
    LessThan_4u_4u LessThan_491 (.cin(1'b0), .a({4'b0000}), .b({delay_counter}), 
            .o(n492));   // insn_decoder.v(531)
    add_4u_4u add_492 (.cin(1'b1), .a({delay_counter}), .b({4'b1110}), 
            .o({n494, n495, n496, n497}));   // insn_decoder.v(531)
    assign n498 = n492 ? n494 : delay_counter[3];   // insn_decoder.v(531)
    assign n499 = n492 ? n495 : delay_counter[2];   // insn_decoder.v(531)
    assign n500 = n492 ? n496 : delay_counter[1];   // insn_decoder.v(531)
    assign n501 = n492 ? n497 : delay_counter[0];   // insn_decoder.v(531)
    nor (n502, n498, n499, n500, n501) ;   // insn_decoder.v(533)
    assign n503 = n502 ? 1'b0 : n39;   // insn_decoder.v(533)
    assign n504 = n502 ? 1'b0 : n40;   // insn_decoder.v(533)
    assign n505 = n502 ? 1'b0 : n41;   // insn_decoder.v(533)
    assign n506 = n502 ? 1'b0 : n42;   // insn_decoder.v(533)
    assign n507 = n502 ? 1'b0 : n43;   // insn_decoder.v(533)
    assign n508 = n502 ? 1'b0 : n44;   // insn_decoder.v(533)
    assign n509 = n502 ? 1'b0 : n45;   // insn_decoder.v(533)
    assign n510 = n502 ? 1'b0 : n46;   // insn_decoder.v(533)
    not (n511, hazard) ;   // insn_decoder.v(540)
    assign n512 = n511 ? old_pcincr_hz : n47;   // insn_decoder.v(540)
    assign n513 = n511 ? old_pass_hz : n48;   // insn_decoder.v(540)
    assign n514 = n511 ? 1'b1 : n49;   // insn_decoder.v(540)
    assign n515 = n511 ? old_fetch_hz : fetch;   // insn_decoder.v(540)
    assign n516 = n511 ? old_state1_hz[7] : n39;   // insn_decoder.v(540)
    assign n517 = n511 ? old_state1_hz[6] : n40;   // insn_decoder.v(540)
    assign n518 = n511 ? old_state1_hz[5] : n41;   // insn_decoder.v(540)
    assign n519 = n511 ? old_state1_hz[4] : n42;   // insn_decoder.v(540)
    assign n520 = n511 ? old_state1_hz[3] : n43;   // insn_decoder.v(540)
    assign n521 = n511 ? old_state1_hz[2] : n44;   // insn_decoder.v(540)
    assign n522 = n511 ? old_state1_hz[1] : n45;   // insn_decoder.v(540)
    assign n523 = n511 ? old_state1_hz[0] : n46;   // insn_decoder.v(540)
    nor (n524, state1[7], state1[6], state1[5], state1[4], state1[3], 
        state1[2], state1[1], state1[0]) ;   // insn_decoder.v(200)
    not (n525, state1[0]) ;   // insn_decoder.v(207)
    nor (n526, state1[7], state1[6], state1[5], state1[4], state1[3], 
        state1[2], state1[1], n525) ;   // insn_decoder.v(207)
    not (n527, state1[1]) ;   // insn_decoder.v(214)
    nor (n528, state1[7], state1[6], state1[5], state1[4], state1[3], 
        state1[2], n527, state1[0]) ;   // insn_decoder.v(214)
    nor (n531, state1[7], state1[6], state1[5], state1[4], state1[3], 
        state1[2], n527, n525) ;   // insn_decoder.v(221)
    not (n532, state1[2]) ;   // insn_decoder.v(228)
    nor (n533, state1[7], state1[6], state1[5], state1[4], state1[3], 
        n532, state1[1], state1[0]) ;   // insn_decoder.v(228)
    nor (n536, state1[7], state1[6], state1[5], state1[4], state1[3], 
        n532, state1[1], n525) ;   // insn_decoder.v(235)
    nor (n539, state1[7], state1[6], state1[5], state1[4], state1[3], 
        n532, n527, state1[0]) ;   // insn_decoder.v(243)
    nor (n546, state1[7], state1[6], state1[5], state1[4], state1[3], 
        n532, n527, n525) ;   // insn_decoder.v(258)
    not (n547, state1[3]) ;   // insn_decoder.v(265)
    nor (n548, state1[7], state1[6], state1[5], state1[4], n547, 
        state1[2], state1[1], state1[0]) ;   // insn_decoder.v(265)
    nor (n551, state1[7], state1[6], state1[5], state1[4], n547, 
        state1[2], state1[1], n525) ;   // insn_decoder.v(272)
    nor (n554, state1[7], state1[6], state1[5], state1[4], n547, 
        state1[2], n527, state1[0]) ;   // insn_decoder.v(279)
    nor (n558, state1[7], state1[6], state1[5], state1[4], n547, 
        state1[2], n527, n525) ;   // insn_decoder.v(286)
    nor (n561, state1[7], state1[6], state1[5], state1[4], n547, 
        n532, state1[1], state1[0]) ;   // insn_decoder.v(293)
    nor (n565, state1[7], state1[6], state1[5], state1[4], n547, 
        n532, state1[1], n525) ;   // insn_decoder.v(301)
    nor (n569, state1[7], state1[6], state1[5], state1[4], n547, 
        n532, n527, state1[0]) ;   // insn_decoder.v(308)
    nor (n574, state1[7], state1[6], state1[5], state1[4], n547, 
        n532, n527, n525) ;   // insn_decoder.v(315)
    not (n575, state1[4]) ;   // insn_decoder.v(322)
    nor (n576, state1[7], state1[6], state1[5], n575, state1[3], 
        state1[2], state1[1], state1[0]) ;   // insn_decoder.v(322)
    nor (n579, state1[7], state1[6], state1[5], n575, state1[3], 
        state1[2], state1[1], n525) ;   // insn_decoder.v(329)
    nor (n582, state1[7], state1[6], state1[5], n575, state1[3], 
        state1[2], n527, state1[0]) ;   // insn_decoder.v(337)
    nor (n586, state1[7], state1[6], state1[5], n575, state1[3], 
        state1[2], n527, n525) ;   // insn_decoder.v(345)
    nor (n589, state1[7], state1[6], state1[5], n575, state1[3], 
        n532, state1[1], state1[0]) ;   // insn_decoder.v(354)
    nor (n593, state1[7], state1[6], state1[5], n575, state1[3], 
        n532, state1[1], n525) ;   // insn_decoder.v(363)
    nor (n597, state1[7], state1[6], state1[5], n575, state1[3], 
        n532, n527, state1[0]) ;   // insn_decoder.v(370)
    nor (n602, state1[7], state1[6], state1[5], n575, state1[3], 
        n532, n527, n525) ;   // insn_decoder.v(377)
    nor (n605, state1[7], state1[6], state1[5], n575, n547, state1[2], 
        state1[1], state1[0]) ;   // insn_decoder.v(385)
    nor (n609, state1[7], state1[6], state1[5], n575, n547, state1[2], 
        state1[1], n525) ;   // insn_decoder.v(398)
    nor (n613, state1[7], state1[6], state1[5], n575, n547, state1[2], 
        n527, state1[0]) ;   // insn_decoder.v(411)
    nor (n618, state1[7], state1[6], state1[5], n575, n547, state1[2], 
        n527, n525) ;   // insn_decoder.v(432)
    nor (n622, state1[7], state1[6], state1[5], n575, n547, n532, 
        state1[1], state1[0]) ;   // insn_decoder.v(445)
    nor (n627, state1[7], state1[6], state1[5], n575, n547, n532, 
        state1[1], n525) ;   // insn_decoder.v(454)
    nor (n632, state1[7], state1[6], state1[5], n575, n547, n532, 
        n527, state1[0]) ;   // insn_decoder.v(472)
    nor (n638, state1[7], state1[6], state1[5], n575, n547, n532, 
        n527, n525) ;   // insn_decoder.v(481)
    not (n639, state1[5]) ;   // insn_decoder.v(495)
    nor (n640, state1[7], state1[6], n639, state1[4], state1[3], 
        state1[2], state1[1], state1[0]) ;   // insn_decoder.v(495)
    nor (n643, state1[7], state1[6], n639, state1[4], state1[3], 
        state1[2], state1[1], n525) ;   // insn_decoder.v(503)
    not (n644, state1[7]) ;   // insn_decoder.v(519)
    nor (n1316, n644, state1[6], state1[5], state1[4], state1[3], 
        state1[2], state1[1], state1[0]) ;   // insn_decoder.v(519)
    nor (n1342, n644, state1[6], state1[5], state1[4], state1[3], 
        state1[2], state1[1], n525) ;   // insn_decoder.v(525)
    nor (n651, n644, state1[6], state1[5], state1[4], state1[3], 
        state1[2], n527, state1[0]) ;   // insn_decoder.v(529)
    nor (n655, n644, state1[6], state1[5], state1[4], state1[3], 
        state1[2], n527, n525) ;   // insn_decoder.v(538)
    not (n656, n524) ;   // insn_decoder.v(198)
    and (n657, n526, n656) ;   // insn_decoder.v(198)
    or (n658, n524, n526) ;   // insn_decoder.v(198)
    not (n659, n658) ;   // insn_decoder.v(198)
    and (n660, n528, n659) ;   // insn_decoder.v(198)
    or (n661, n658, n528) ;   // insn_decoder.v(198)
    not (n662, n661) ;   // insn_decoder.v(198)
    and (n663, n531, n662) ;   // insn_decoder.v(198)
    or (n664, n661, n531) ;   // insn_decoder.v(198)
    not (n665, n664) ;   // insn_decoder.v(198)
    and (n666, n533, n665) ;   // insn_decoder.v(198)
    or (n667, n664, n533) ;   // insn_decoder.v(198)
    not (n668, n667) ;   // insn_decoder.v(198)
    and (n669, n536, n668) ;   // insn_decoder.v(198)
    or (n670, n667, n536) ;   // insn_decoder.v(198)
    not (n671, n670) ;   // insn_decoder.v(198)
    and (n672, n539, n671) ;   // insn_decoder.v(198)
    or (n673, n670, n539) ;   // insn_decoder.v(198)
    not (n674, n673) ;   // insn_decoder.v(198)
    and (n675, n539, n674) ;   // insn_decoder.v(198)
    or (n676, n673, n539) ;   // insn_decoder.v(198)
    not (n677, n676) ;   // insn_decoder.v(198)
    and (n678, n546, n677) ;   // insn_decoder.v(198)
    or (n679, n676, n546) ;   // insn_decoder.v(198)
    not (n680, n679) ;   // insn_decoder.v(198)
    and (n681, n548, n680) ;   // insn_decoder.v(198)
    or (n682, n679, n548) ;   // insn_decoder.v(198)
    not (n683, n682) ;   // insn_decoder.v(198)
    and (n684, n551, n683) ;   // insn_decoder.v(198)
    or (n685, n682, n551) ;   // insn_decoder.v(198)
    not (n686, n685) ;   // insn_decoder.v(198)
    and (n687, n554, n686) ;   // insn_decoder.v(198)
    or (n688, n685, n554) ;   // insn_decoder.v(198)
    not (n689, n688) ;   // insn_decoder.v(198)
    and (n690, n558, n689) ;   // insn_decoder.v(198)
    or (n691, n688, n558) ;   // insn_decoder.v(198)
    not (n692, n691) ;   // insn_decoder.v(198)
    and (n693, n561, n692) ;   // insn_decoder.v(198)
    or (n694, n691, n561) ;   // insn_decoder.v(198)
    not (n695, n694) ;   // insn_decoder.v(198)
    and (n696, n565, n695) ;   // insn_decoder.v(198)
    or (n697, n694, n565) ;   // insn_decoder.v(198)
    not (n698, n697) ;   // insn_decoder.v(198)
    and (n699, n569, n698) ;   // insn_decoder.v(198)
    or (n700, n697, n569) ;   // insn_decoder.v(198)
    not (n701, n700) ;   // insn_decoder.v(198)
    and (n702, n574, n701) ;   // insn_decoder.v(198)
    or (n703, n700, n574) ;   // insn_decoder.v(198)
    not (n704, n703) ;   // insn_decoder.v(198)
    and (n705, n576, n704) ;   // insn_decoder.v(198)
    or (n706, n703, n576) ;   // insn_decoder.v(198)
    not (n707, n706) ;   // insn_decoder.v(198)
    and (n708, n579, n707) ;   // insn_decoder.v(198)
    or (n709, n706, n579) ;   // insn_decoder.v(198)
    not (n710, n709) ;   // insn_decoder.v(198)
    and (n711, n582, n710) ;   // insn_decoder.v(198)
    or (n712, n709, n582) ;   // insn_decoder.v(198)
    not (n713, n712) ;   // insn_decoder.v(198)
    and (n714, n586, n713) ;   // insn_decoder.v(198)
    or (n715, n712, n586) ;   // insn_decoder.v(198)
    not (n716, n715) ;   // insn_decoder.v(198)
    and (n717, n589, n716) ;   // insn_decoder.v(198)
    or (n718, n715, n589) ;   // insn_decoder.v(198)
    not (n719, n718) ;   // insn_decoder.v(198)
    and (n720, n593, n719) ;   // insn_decoder.v(198)
    or (n721, n718, n593) ;   // insn_decoder.v(198)
    not (n722, n721) ;   // insn_decoder.v(198)
    and (n723, n597, n722) ;   // insn_decoder.v(198)
    or (n724, n721, n597) ;   // insn_decoder.v(198)
    not (n725, n724) ;   // insn_decoder.v(198)
    and (n726, n602, n725) ;   // insn_decoder.v(198)
    or (n727, n724, n602) ;   // insn_decoder.v(198)
    not (n728, n727) ;   // insn_decoder.v(198)
    and (n729, n605, n728) ;   // insn_decoder.v(198)
    or (n730, n727, n605) ;   // insn_decoder.v(198)
    not (n731, n730) ;   // insn_decoder.v(198)
    and (n732, n609, n731) ;   // insn_decoder.v(198)
    or (n733, n730, n609) ;   // insn_decoder.v(198)
    not (n734, n733) ;   // insn_decoder.v(198)
    and (n735, n613, n734) ;   // insn_decoder.v(198)
    or (n736, n733, n613) ;   // insn_decoder.v(198)
    not (n737, n736) ;   // insn_decoder.v(198)
    and (n738, n618, n737) ;   // insn_decoder.v(198)
    or (n739, n736, n618) ;   // insn_decoder.v(198)
    not (n740, n739) ;   // insn_decoder.v(198)
    and (n741, n622, n740) ;   // insn_decoder.v(198)
    or (n742, n739, n622) ;   // insn_decoder.v(198)
    not (n743, n742) ;   // insn_decoder.v(198)
    and (n744, n627, n743) ;   // insn_decoder.v(198)
    or (n745, n742, n627) ;   // insn_decoder.v(198)
    not (n746, n745) ;   // insn_decoder.v(198)
    and (n747, n632, n746) ;   // insn_decoder.v(198)
    or (n748, n745, n632) ;   // insn_decoder.v(198)
    not (n749, n748) ;   // insn_decoder.v(198)
    and (n750, n638, n749) ;   // insn_decoder.v(198)
    or (n751, n748, n638) ;   // insn_decoder.v(198)
    not (n752, n751) ;   // insn_decoder.v(198)
    and (n753, n640, n752) ;   // insn_decoder.v(198)
    or (n754, n751, n640) ;   // insn_decoder.v(198)
    not (n755, n754) ;   // insn_decoder.v(198)
    and (n756, n643, n755) ;   // insn_decoder.v(198)
    or (n757, n754, n643) ;   // insn_decoder.v(198)
    not (n758, n757) ;   // insn_decoder.v(198)
    and (n759, n1316, n758) ;   // insn_decoder.v(198)
    or (n760, n757, n1316) ;   // insn_decoder.v(198)
    not (n761, n760) ;   // insn_decoder.v(198)
    and (n762, n1342, n761) ;   // insn_decoder.v(198)
    or (n763, n760, n1342) ;   // insn_decoder.v(198)
    not (n764, n763) ;   // insn_decoder.v(198)
    and (n765, n651, n764) ;   // insn_decoder.v(198)
    or (n766, n763, n651) ;   // insn_decoder.v(198)
    not (n767, n766) ;   // insn_decoder.v(198)
    and (n768, n655, n767) ;   // insn_decoder.v(198)
    or (n769, n766, n655) ;   // insn_decoder.v(198)
    not (n770, n769) ;   // insn_decoder.v(198)
    or (n771, n759, n762, n765, n768, n770) ;   // insn_decoder.v(198)
    assign n772 = n771 ? e_alu_op[7] : 1'b0;   // insn_decoder.v(198)
    assign n774 = n771 ? e_alu_op[6] : 1'b0;   // insn_decoder.v(198)
    assign n776 = n771 ? e_alu_op[5] : 1'b0;   // insn_decoder.v(198)
    or (n777, n524, n657, n663, n666, n669, n672, n678, n681, 
        n684, n687, n690, n693, n696, n699, n702, n705, n708, 
        n711, n714, n717, n720, n723, n726, n729, n732, n735, 
        n738, n741, n744, n747, n750, n753, n756) ;   // insn_decoder.v(198)
    or (n778, n660, n675) ;   // insn_decoder.v(198)
    Select_3 Select_775 (.sel({n777, n778, n771}), .data({2'b01, e_alu_op[4]}), 
            .o(n780));   // insn_decoder.v(198)
    or (n781, n524, n660, n675, n678, n681, n684, n696, n699, 
            n702, n705, n708, n711, n714, n717, n720, n723, 
            n729, n732, n735, n738, n741, n744, n747, n750, 
            n753, n756) ;   // insn_decoder.v(198)
    or (n782, n657, n663, n666, n669, n672, n687, n690, n693, 
            n726) ;   // insn_decoder.v(198)
    Select_3 Select_779 (.sel({n781, n782, n771}), .data({2'b01, e_alu_op[3]}), 
            .o(n784));   // insn_decoder.v(198)
    or (n785, n524, n660, n669, n675, n687, n690, n693, n696, 
            n699, n711, n714, n717, n720, n723, n729, n732, 
            n735, n738, n741, n744, n747, n750, n753, n756) ;   // insn_decoder.v(198)
    or (n786, n657, n663, n666, n672, n678, n681, n684, n702, 
            n705, n708, n726) ;   // insn_decoder.v(198)
    Select_3 Select_783 (.sel({n785, n786, n771}), .data({2'b01, e_alu_op[2]}), 
            .o(n788));   // insn_decoder.v(198)
    or (n789, n524, n657, n660, n663, n675, n681, n687, n690, 
            n696, n702, n705, n708, n714, n723, n726, n729, 
            n732, n735, n738, n741, n744, n747, n750, n753, 
            n756) ;   // insn_decoder.v(198)
    or (n790, n666, n669, n672, n678, n684, n693, n699, n711, 
            n717, n720) ;   // insn_decoder.v(198)
    Select_3 Select_787 (.sel({n789, n790, n771}), .data({2'b01, e_alu_op[1]}), 
            .o(n792));   // insn_decoder.v(198)
    or (n793, n524, n660, n663, n672, n678, n687, n693, n699, 
            n702, n705, n708, n717, n720, n726, n729, n735, 
            n738, n741, n744, n747, n750, n753, n756) ;   // insn_decoder.v(198)
    or (n794, n657, n666, n669, n675, n681, n684, n690, n696, 
            n711, n714, n723, n732) ;   // insn_decoder.v(198)
    Select_3 Select_791 (.sel({n793, n794, n771}), .data({2'b01, e_alu_op[0]}), 
            .o(n796));   // insn_decoder.v(198)
    or (n797, n657, n660, n663, n666, n669, n672, n675, n678, 
            n681, n684, n687, n690, n693, n696, n699, n702, 
            n705, n708, n711, n714, n717, n720, n723, n726, 
            n729, n732, n735, n738, n741, n744, n747, n750, 
            n753, n756) ;   // insn_decoder.v(198)
    Select_3 Select_794 (.sel({n524, n797, n771}), .data({1'b0, cond[3], 
            e_cond[3]}), .o(n799));   // insn_decoder.v(198)
    Select_3 Select_797 (.sel({n524, n797, n771}), .data({1'b0, cond[2], 
            e_cond[2]}), .o(n802));   // insn_decoder.v(198)
    Select_3 Select_800 (.sel({n524, n797, n771}), .data({1'b0, cond[1], 
            e_cond[1]}), .o(n805));   // insn_decoder.v(198)
    Select_3 Select_803 (.sel({n524, n797, n771}), .data({1'b0, cond[0], 
            e_cond[0]}), .o(n808));   // insn_decoder.v(198)
    or (n809, n524, n729, n732, n735, n738, n741, n744, n747, 
            n750, n753, n756) ;   // insn_decoder.v(198)
    or (n810, n657, n660, n663, n666, n669, n672, n675, n678, 
            n681, n684, n687, n690, n693, n696, n699, n702, 
            n705, n708, n711, n714, n717, n720, n723, n726) ;   // insn_decoder.v(198)
    Select_3 Select_807 (.sel({n809, n810, n771}), .data({2'b01, e_write_flags[3]}), 
            .o(n812));   // insn_decoder.v(198)
    Select_3 Select_811 (.sel({n809, n810, n771}), .data({2'b01, e_write_flags[2]}), 
            .o(n816));   // insn_decoder.v(198)
    Select_3 Select_815 (.sel({n809, n810, n771}), .data({2'b01, e_write_flags[1]}), 
            .o(n820));   // insn_decoder.v(198)
    Select_3 Select_819 (.sel({n809, n810, n771}), .data({2'b01, e_write_flags[0]}), 
            .o(n824));   // insn_decoder.v(198)
    Select_3 Select_822 (.sel({n524, n797, n771}), .data({2'b01, e_is_cond}), 
            .o(n827));   // insn_decoder.v(198)
    or (n828, n524, n657, n660, n663, n666, n669, n672, n675, 
            n678, n681, n684, n687, n690, n693, n696, n699, 
            n702, n705, n708, n711, n714, n717, n720, n723, 
            n726, n729, n732, n735, n738, n741, n744, n750, 
            n753, n756) ;   // insn_decoder.v(198)
    Select_3 Select_825 (.sel({n828, n747, n771}), .data({2'b01, m_r1_op[3]}), 
            .o(n830));   // insn_decoder.v(198)
    assign n832 = n771 ? m_r1_op[2] : 1'b0;   // insn_decoder.v(198)
    or (n833, n524, n657, n660, n663, n666, n669, n672, n675, 
        n678, n681, n684, n687, n690, n693, n696, n699, n702, 
        n705, n708, n711, n714, n717, n720, n723, n726, n729, 
        n732, n735, n738, n744, n747, n750, n753, n756) ;   // insn_decoder.v(198)
    Select_3 Select_830 (.sel({n833, n741, n771}), .data({2'b01, m_r1_op[1]}), 
            .o(n835));   // insn_decoder.v(198)
    or (n836, n524, n741, n747) ;   // insn_decoder.v(198)
    or (n837, n657, n660, n663, n666, n669, n672, n675, n678, 
            n681, n684, n687, n690, n693, n696, n699, n702, 
            n705, n708, n711, n714, n717, n720, n723, n726, 
            n729, n732, n735, n738, n744, n750, n753, n756) ;   // insn_decoder.v(198)
    Select_3 Select_834 (.sel({n836, n837, n771}), .data({2'b01, m_r1_op[0]}), 
            .o(n839));   // insn_decoder.v(198)
    or (n840, n524, n657, n660, n663, n666, n669, n672, n675, 
            n678, n681, n684, n687, n690, n693, n696, n699, 
            n702, n705, n708, n711, n714, n717, n720, n723, 
            n726, n729, n732, n735, n738, n741, n744, n747, 
            n753, n756) ;   // insn_decoder.v(198)
    Select_3 Select_837 (.sel({n840, n750, n771}), .data({2'b01, m_r2_op[3]}), 
            .o(n842));   // insn_decoder.v(198)
    or (n843, n524, n657, n660, n663, n666, n669, n672, n675, 
            n678, n681, n684, n687, n690, n693, n696, n699, 
            n702, n705, n708, n711, n714, n717, n720, n723, 
            n726, n729, n732, n735, n738, n741, n747, n750, 
            n753, n756) ;   // insn_decoder.v(198)
    Select_3 Select_840 (.sel({n843, n744, n771}), .data({2'b01, m_r2_op[2]}), 
            .o(n845));   // insn_decoder.v(198)
    Select_3 Select_843 (.sel({n840, n750, n771}), .data({2'b01, m_r2_op[1]}), 
            .o(n848));   // insn_decoder.v(198)
    Select_3 Select_846 (.sel({n524, n797, n771}), .data({2'b01, m_r2_op[0]}), 
            .o(n851));   // insn_decoder.v(198)
    assign n853 = n771 ? r_op[3] : 1'b0;   // insn_decoder.v(198)
    or (n854, n524, n657, n660, n663, n666, n669, n672, n675, 
        n678, n681, n684, n687, n690, n693, n696, n699, n702, 
        n711, n714, n717, n720, n723, n726, n729, n732, n738, 
        n741, n744, n747, n750, n753) ;   // insn_decoder.v(198)
    or (n855, n705, n708, n735, n756) ;   // insn_decoder.v(198)
    Select_3 Select_852 (.sel({n854, n855, n771}), .data({2'b01, r_op[2]}), 
            .o(n857));   // insn_decoder.v(198)
    or (n858, n524, n657, n660, n663, n666, n669, n672, n675, 
            n678, n681, n684, n687, n690, n693, n696, n699, 
            n702, n705, n711, n714, n717, n720, n723, n726, 
            n729, n732, n738, n741, n744, n747, n750, n753) ;   // insn_decoder.v(198)
    or (n859, n708, n735, n756) ;   // insn_decoder.v(198)
    Select_3 Select_856 (.sel({n858, n859, n771}), .data({2'b01, r_op[1]}), 
            .o(n861));   // insn_decoder.v(198)
    or (n862, n524, n705, n720, n723, n726, n744, n750) ;   // insn_decoder.v(198)
    or (n863, n657, n660, n663, n666, n669, n672, n675, n678, 
            n681, n684, n687, n690, n693, n696, n699, n702, 
            n708, n711, n714, n717, n729, n732, n735, n738, 
            n741, n747, n753, n756) ;   // insn_decoder.v(198)
    Select_3 Select_860 (.sel({n862, n863, n771}), .data({2'b01, r_op[0]}), 
            .o(n865));   // insn_decoder.v(198)
    or (n866, n524, n669, n711, n714, n717, n729, n738, n741, 
            n747, n753) ;   // insn_decoder.v(198)
    or (n867, n657, n660, n663, n666, n672, n675, n678, n681, 
            n684, n687, n690, n693, n696, n699, n702, n705, 
            n708, n720, n723, n726, n732, n735, n744, n750, 
            n756) ;   // insn_decoder.v(198)
    Select_3 Select_864 (.sel({n866, n867, n771}), .data({2'b01, r_read[1]}), 
            .o(n869));   // insn_decoder.v(198)
    Select_3 Select_867 (.sel({n524, n797, n771}), .data({2'b01, r_read[0]}), 
            .o(n872));   // insn_decoder.v(198)
    assign n874 = n771 ? r_to_mem[1] : 1'b0;   // insn_decoder.v(198)
    or (n875, n524, n657, n660, n663, n666, n669, n672, n675, 
        n678, n681, n684, n687, n690, n693, n696, n699, n702, 
        n705, n708, n711, n714, n717, n720, n723, n726, n729, 
        n732, n735, n738, n753, n756) ;   // insn_decoder.v(198)
    or (n876, n741, n744, n747, n750) ;   // insn_decoder.v(198)
    Select_3 Select_873 (.sel({n875, n876, n771}), .data({2'b01, r_to_mem[0]}), 
            .o(n878));   // insn_decoder.v(198)
    or (n879, n524, n720, n723, n726, n744, n750, n759, n762, 
            n765, n768, n770) ;   // insn_decoder.v(198)
    or (n880, n657, n660, n663, n666, n669, n672, n675, n678, 
            n681, n684, n687, n690, n693, n696, n699, n702, 
            n705, n708, n711, n714, n717, n741, n747, n753, 
            n756) ;   // insn_decoder.v(198)
    or (n881, n729, n732, n735, n738) ;   // insn_decoder.v(198)
    Select_3 Select_877 (.sel({n879, n880, n881}), .data({r_a1[4], reg_c_addr[4], 
            1'b1}), .o(n882));   // insn_decoder.v(198)
    Select_3 Select_881 (.sel({n879, n880, n881}), .data({r_a1[3], reg_c_addr[3], 
            1'b1}), .o(n886));   // insn_decoder.v(198)
    Select_3 Select_885 (.sel({n879, n880, n881}), .data({r_a1[2], reg_c_addr[2], 
            1'b1}), .o(n890));   // insn_decoder.v(198)
    Select_3 Select_889 (.sel({n879, n880, n881}), .data({r_a1[1], reg_c_addr[1], 
            1'b1}), .o(n894));   // insn_decoder.v(198)
    Select_3 Select_893 (.sel({n879, n880, n881}), .data({r_a1[0], reg_c_addr[0], 
            1'b1}), .o(n898));   // insn_decoder.v(198)
    or (n899, n524, n759, n762, n765, n768, n770) ;   // insn_decoder.v(198)
    or (n900, n657, n660, n663, n666, n669, n672, n675, n678, 
            n681, n684, n687, n690, n693, n696, n699, n702, 
            n705, n708, n711, n714, n717, n720, n723, n726, 
            n729, n735, n741, n744, n747, n750, n753, n756) ;   // insn_decoder.v(198)
    or (n901, n732, n738) ;   // insn_decoder.v(198)
    Select_3 Select_897 (.sel({n899, n900, n901}), .data({r_r1_addr[4], 
            reg_a_addr[4], 1'b1}), .o(n902));   // insn_decoder.v(198)
    Select_3 Select_901 (.sel({n899, n900, n901}), .data({r_r1_addr[3], 
            reg_a_addr[3], 1'b1}), .o(n906));   // insn_decoder.v(198)
    Select_3 Select_905 (.sel({n899, n900, n901}), .data({r_r1_addr[2], 
            reg_a_addr[2], 1'b1}), .o(n910));   // insn_decoder.v(198)
    Select_4 Select_908 (.sel({n899, n900, n732, n738}), .data({r_r1_addr[1], 
            reg_a_addr[1], 2'b10}), .o(n913));   // insn_decoder.v(198)
    Select_3 Select_912 (.sel({n899, n900, n901}), .data({r_r1_addr[0], 
            reg_a_addr[0], 1'b1}), .o(n917));   // insn_decoder.v(198)
    or (n918, n524, n669, n711, n714, n717, n729, n738, n741, 
            n747, n753, n759, n762, n765, n768, n770) ;   // insn_decoder.v(198)
    or (n919, n657, n660, n663, n666, n672, n675, n678, n681, 
            n684, n687, n690, n693, n696, n699, n702, n705, 
            n708, n720, n723, n726, n744, n750, n756) ;   // insn_decoder.v(198)
    Select_4 Select_915 (.sel({n918, n919, n732, n735}), .data({r_r2_addr[4], 
            reg_b_addr[4], reg_a_addr[4], 1'b1}), .o(n920));   // insn_decoder.v(198)
    Select_4 Select_918 (.sel({n918, n919, n732, n735}), .data({r_r2_addr[3], 
            reg_b_addr[3], reg_a_addr[3], 1'b1}), .o(n923));   // insn_decoder.v(198)
    Select_4 Select_921 (.sel({n918, n919, n732, n735}), .data({r_r2_addr[2], 
            reg_b_addr[2], reg_a_addr[2], 1'b1}), .o(n926));   // insn_decoder.v(198)
    Select_4 Select_924 (.sel({n918, n919, n732, n735}), .data({r_r2_addr[1], 
            reg_b_addr[1], reg_a_addr[1], 1'b1}), .o(n929));   // insn_decoder.v(198)
    Select_4 Select_927 (.sel({n918, n919, n732, n735}), .data({r_r2_addr[0], 
            reg_b_addr[0], reg_a_addr[0], 1'b1}), .o(n932));   // insn_decoder.v(198)
    or (n933, n524, n657, n660, n663, n666, n669, n672, n675, 
            n678, n681, n684, n687, n690, n693, n696, n699, 
            n702, n705, n711, n714, n717, n720, n723, n726, 
            n729, n732, n735, n753, n759, n762, n765, n768, 
            n770) ;   // insn_decoder.v(198)
    or (n934, n708, n738, n756) ;   // insn_decoder.v(198)
    Select_3 Select_931 (.sel({n933, n934, n876}), .data({n36, 2'b01}), 
            .o(n936));   // insn_decoder.v(198)
    assign n939 = n934 ? 1'b0 : n37;   // insn_decoder.v(198)
    or (n941, n669, n708, n711, n714, n717, n729, n732, n735, 
        n738, n741, n744, n747, n750, n753, n756) ;   // insn_decoder.v(198)
    assign n942 = n941 ? 1'b0 : n38;   // insn_decoder.v(198)
    or (n943, n524, n657, n660, n663, n666, n669, n672, n675, 
        n678, n681, n684, n687, n690, n693, n696, n699, n702, 
        n705, n711, n714, n717, n720, n723, n726, n729, n732, 
        n738, n741, n744, n747, n750, n753, n759, n762, n765, 
        n768, n770) ;   // insn_decoder.v(198)
    or (n944, n708, n756) ;   // insn_decoder.v(198)
    Select_3 Select_940 (.sel({n943, n944, n735}), .data({r_a2[4], reg_d_addr[4], 
            1'b1}), .o(n945));   // insn_decoder.v(198)
    Select_3 Select_943 (.sel({n943, n944, n735}), .data({r_a2[3], reg_d_addr[3], 
            1'b1}), .o(n948));   // insn_decoder.v(198)
    Select_3 Select_946 (.sel({n943, n944, n735}), .data({r_a2[2], reg_d_addr[2], 
            1'b1}), .o(n951));   // insn_decoder.v(198)
    Select_3 Select_949 (.sel({n943, n944, n735}), .data({r_a2[1], reg_d_addr[1], 
            1'b0}), .o(n954));   // insn_decoder.v(198)
    Select_3 Select_952 (.sel({n943, n944, n735}), .data({r_a2[0], reg_d_addr[0], 
            1'b1}), .o(n957));   // insn_decoder.v(198)
    or (n958, n524, n657, n660, n663, n666, n669, n672, n675, 
            n678, n681, n684, n687, n690, n693, n696, n699, 
            n702, n705, n708, n711, n720, n723, n726, n729, 
            n732, n735, n738, n741, n744, n747, n750, n753, 
            n756, n765, n768, n770) ;   // insn_decoder.v(198)
    or (n959, n714, n717) ;   // insn_decoder.v(198)
    Select_4 Select_955 (.sel({n958, n959, n759, n762}), .data({e_b[31], 
            1'b0, n261, n428}), .o(n960));   // insn_decoder.v(198)
    Select_4 Select_958 (.sel({n958, n959, n759, n762}), .data({e_b[30], 
            1'b0, n262, n429}), .o(n963));   // insn_decoder.v(198)
    Select_4 Select_961 (.sel({n958, n959, n759, n762}), .data({e_b[29], 
            1'b0, n263, n430}), .o(n966));   // insn_decoder.v(198)
    Select_4 Select_964 (.sel({n958, n959, n759, n762}), .data({e_b[28], 
            1'b0, n264, n431}), .o(n969));   // insn_decoder.v(198)
    Select_4 Select_967 (.sel({n958, n959, n759, n762}), .data({e_b[27], 
            1'b0, n265, n432}), .o(n972));   // insn_decoder.v(198)
    Select_4 Select_970 (.sel({n958, n959, n759, n762}), .data({e_b[26], 
            1'b0, n266, n433}), .o(n975));   // insn_decoder.v(198)
    Select_4 Select_973 (.sel({n958, n959, n759, n762}), .data({e_b[25], 
            1'b0, n267, n434}), .o(n978));   // insn_decoder.v(198)
    Select_4 Select_976 (.sel({n958, n959, n759, n762}), .data({e_b[24], 
            1'b0, n268, n435}), .o(n981));   // insn_decoder.v(198)
    Select_4 Select_979 (.sel({n958, n959, n759, n762}), .data({e_b[23], 
            1'b0, n269, n436}), .o(n984));   // insn_decoder.v(198)
    Select_4 Select_982 (.sel({n958, n959, n759, n762}), .data({e_b[22], 
            1'b0, n270, n437}), .o(n987));   // insn_decoder.v(198)
    Select_4 Select_985 (.sel({n958, n959, n759, n762}), .data({e_b[21], 
            1'b0, n271, n438}), .o(n990));   // insn_decoder.v(198)
    Select_4 Select_988 (.sel({n958, n959, n759, n762}), .data({e_b[20], 
            1'b0, n272, n439}), .o(n993));   // insn_decoder.v(198)
    Select_4 Select_991 (.sel({n958, n959, n759, n762}), .data({e_b[19], 
            1'b0, n273, n440}), .o(n996));   // insn_decoder.v(198)
    Select_4 Select_994 (.sel({n958, n959, n759, n762}), .data({e_b[18], 
            1'b0, n274, n441}), .o(n999));   // insn_decoder.v(198)
    Select_4 Select_997 (.sel({n958, n959, n759, n762}), .data({e_b[17], 
            1'b0, n275, n442}), .o(n1002));   // insn_decoder.v(198)
    Select_4 Select_1000 (.sel({n958, n959, n759, n762}), .data({e_b[16], 
            1'b0, n276, n443}), .o(n1005));   // insn_decoder.v(198)
    Select_4 Select_1003 (.sel({n958, n959, n759, n762}), .data({e_b[15], 
            1'b0, n277, n444}), .o(n1008));   // insn_decoder.v(198)
    Select_4 Select_1006 (.sel({n958, n959, n759, n762}), .data({e_b[14], 
            1'b0, n278, n445}), .o(n1011));   // insn_decoder.v(198)
    Select_4 Select_1009 (.sel({n958, n959, n759, n762}), .data({e_b[13], 
            1'b0, n279, n446}), .o(n1014));   // insn_decoder.v(198)
    Select_4 Select_1012 (.sel({n958, n959, n759, n762}), .data({e_b[12], 
            1'b0, n280, n447}), .o(n1017));   // insn_decoder.v(198)
    Select_4 Select_1015 (.sel({n958, n959, n759, n762}), .data({e_b[11], 
            1'b0, n281, n448}), .o(n1020));   // insn_decoder.v(198)
    Select_4 Select_1018 (.sel({n958, n959, n759, n762}), .data({e_b[10], 
            1'b0, n282, n449}), .o(n1023));   // insn_decoder.v(198)
    Select_4 Select_1021 (.sel({n958, n959, n759, n762}), .data({e_b[9], 
            1'b0, n283, n450}), .o(n1026));   // insn_decoder.v(198)
    Select_4 Select_1024 (.sel({n958, n959, n759, n762}), .data({e_b[8], 
            1'b0, n284, n451}), .o(n1029));   // insn_decoder.v(198)
    Select_4 Select_1027 (.sel({n958, n959, n759, n762}), .data({e_b[7], 
            1'b0, n285, n452}), .o(n1032));   // insn_decoder.v(198)
    Select_4 Select_1030 (.sel({n958, n959, n759, n762}), .data({e_b[6], 
            1'b0, n286, n453}), .o(n1035));   // insn_decoder.v(198)
    Select_4 Select_1033 (.sel({n958, n959, n759, n762}), .data({e_b[5], 
            1'b0, n287, n454}), .o(n1038));   // insn_decoder.v(198)
    Select_4 Select_1036 (.sel({n958, n959, n759, n762}), .data({e_b[4], 
            1'b0, n288, n455}), .o(n1041));   // insn_decoder.v(198)
    Select_4 Select_1039 (.sel({n958, n959, n759, n762}), .data({e_b[3], 
            1'b0, n289, n456}), .o(n1044));   // insn_decoder.v(198)
    Select_4 Select_1042 (.sel({n958, n959, n759, n762}), .data({e_b[2], 
            1'b0, n290, n457}), .o(n1047));   // insn_decoder.v(198)
    Select_4 Select_1045 (.sel({n958, n959, n759, n762}), .data({e_b[1], 
            1'b0, n291, n458}), .o(n1050));   // insn_decoder.v(198)
    Select_4 Select_1048 (.sel({n958, n959, n759, n762}), .data({e_b[0], 
            1'b1, n292, n459}), .o(n1053));   // insn_decoder.v(198)
    or (n1054, n524, n657, n660, n663, n666, n669, n672, n675, 
            n678, n681, n684, n687, n690, n693, n696, n699, 
            n702, n705, n708, n711, n714, n717, n720, n723, 
            n726, n741, n744, n747, n750, n753, n756, n759, 
            n762) ;   // insn_decoder.v(198)
    Select_5 Select_1051 (.sel({n1054, n881, n765, n768, n770}), .data({fetch, 
            1'b0, n502, n515, 1'b1}), .o(n1056));   // insn_decoder.v(198)
    or (n1057, n524, n657, n660, n663, n666, n669, n672, n675, 
            n678, n681, n684, n687, n690, n693, n696, n699, 
            n702, n705, n708, n711, n714, n717, n720, n723, 
            n726, n741, n744, n747, n750, n753, n756, n759, 
            n762, n770) ;   // insn_decoder.v(198)
    Select_4 Select_1054 (.sel({n1057, n881, n765, n768}), .data({n47, 
            1'b0, n502, n512}), .o(n1059));   // insn_decoder.v(198)
    Select_5 Select_1057 (.sel({n1054, n881, n765, n768, n770}), .data({n39, 
            1'b1, n503, n516, 1'b0}), .o(n1062));   // insn_decoder.v(198)
    or (n1064, n729, n732, n735, n738, n770) ;   // insn_decoder.v(198)
    Select_4 Select_1060 (.sel({n1054, n1064, n765, n768}), .data({n40, 
            1'b0, n504, n517}), .o(n1065));   // insn_decoder.v(198)
    Select_4 Select_1063 (.sel({n1054, n1064, n765, n768}), .data({n41, 
            1'b0, n505, n518}), .o(n1068));   // insn_decoder.v(198)
    Select_4 Select_1066 (.sel({n1054, n1064, n765, n768}), .data({n42, 
            1'b0, n506, n519}), .o(n1071));   // insn_decoder.v(198)
    Select_4 Select_1069 (.sel({n1054, n1064, n765, n768}), .data({n43, 
            1'b0, n507, n520}), .o(n1074));   // insn_decoder.v(198)
    Select_4 Select_1072 (.sel({n1054, n1064, n765, n768}), .data({n44, 
            1'b0, n508, n521}), .o(n1077));   // insn_decoder.v(198)
    Select_5 Select_1075 (.sel({n1054, n881, n765, n768, n770}), .data({n45, 
            1'b1, n509, n522, 1'b0}), .o(n1080));   // insn_decoder.v(198)
    Select_4 Select_1078 (.sel({n1054, n1064, n765, n768}), .data({n46, 
            1'b0, n510, n523}), .o(n1083));   // insn_decoder.v(198)
    or (n1084, n524, n657, n660, n663, n666, n669, n672, n675, 
            n678, n681, n684, n687, n690, n693, n696, n699, 
            n702, n705, n708, n711, n714, n717, n720, n723, 
            n726, n741, n744, n747, n750, n753, n756, n759, 
            n762, n768, n770) ;   // insn_decoder.v(198)
    Select_3 Select_1081 (.sel({n1084, n881, n765}), .data({delay_counter[3], 
            1'b0, n498}), .o(n1086));   // insn_decoder.v(198)
    Select_3 Select_1084 (.sel({n1084, n881, n765}), .data({delay_counter[2], 
            1'b0, n499}), .o(n1089));   // insn_decoder.v(198)
    Select_3 Select_1087 (.sel({n1084, n881, n765}), .data({delay_counter[1], 
            1'b1, n500}), .o(n1092));   // insn_decoder.v(198)
    Select_3 Select_1090 (.sel({n1084, n881, n765}), .data({delay_counter[0], 
            1'b1, n501}), .o(n1095));   // insn_decoder.v(198)
    assign n1097 = n759 ? n293 : e_a[31];   // insn_decoder.v(198)
    assign n1099 = n759 ? n294 : e_a[30];   // insn_decoder.v(198)
    assign n1101 = n759 ? n295 : e_a[29];   // insn_decoder.v(198)
    assign n1103 = n759 ? n296 : e_a[28];   // insn_decoder.v(198)
    assign n1105 = n759 ? n297 : e_a[27];   // insn_decoder.v(198)
    assign n1107 = n759 ? n298 : e_a[26];   // insn_decoder.v(198)
    assign n1109 = n759 ? n299 : e_a[25];   // insn_decoder.v(198)
    assign n1111 = n759 ? n300 : e_a[24];   // insn_decoder.v(198)
    assign n1113 = n759 ? n301 : e_a[23];   // insn_decoder.v(198)
    assign n1115 = n759 ? n302 : e_a[22];   // insn_decoder.v(198)
    assign n1117 = n759 ? n303 : e_a[21];   // insn_decoder.v(198)
    assign n1119 = n759 ? n304 : e_a[20];   // insn_decoder.v(198)
    assign n1121 = n759 ? n305 : e_a[19];   // insn_decoder.v(198)
    assign n1123 = n759 ? n306 : e_a[18];   // insn_decoder.v(198)
    assign n1125 = n759 ? n307 : e_a[17];   // insn_decoder.v(198)
    assign n1127 = n759 ? n308 : e_a[16];   // insn_decoder.v(198)
    assign n1129 = n759 ? n309 : e_a[15];   // insn_decoder.v(198)
    assign n1131 = n759 ? n310 : e_a[14];   // insn_decoder.v(198)
    assign n1133 = n759 ? n311 : e_a[13];   // insn_decoder.v(198)
    assign n1135 = n759 ? n312 : e_a[12];   // insn_decoder.v(198)
    assign n1137 = n759 ? n313 : e_a[11];   // insn_decoder.v(198)
    assign n1139 = n759 ? n314 : e_a[10];   // insn_decoder.v(198)
    assign n1141 = n759 ? n315 : e_a[9];   // insn_decoder.v(198)
    assign n1143 = n759 ? n316 : e_a[8];   // insn_decoder.v(198)
    assign n1145 = n759 ? n317 : e_a[7];   // insn_decoder.v(198)
    assign n1147 = n759 ? n318 : e_a[6];   // insn_decoder.v(198)
    assign n1149 = n759 ? n319 : e_a[5];   // insn_decoder.v(198)
    assign n1151 = n759 ? n320 : e_a[4];   // insn_decoder.v(198)
    assign n1153 = n759 ? n321 : e_a[3];   // insn_decoder.v(198)
    assign n1155 = n759 ? n322 : e_a[2];   // insn_decoder.v(198)
    assign n1157 = n759 ? n323 : e_a[1];   // insn_decoder.v(198)
    assign n1159 = n759 ? n324 : e_a[0];   // insn_decoder.v(198)
    assign n1161 = n759 ? n325 : m_a1[31];   // insn_decoder.v(198)
    assign n1163 = n759 ? n326 : m_a1[30];   // insn_decoder.v(198)
    assign n1165 = n759 ? n327 : m_a1[29];   // insn_decoder.v(198)
    assign n1167 = n759 ? n328 : m_a1[28];   // insn_decoder.v(198)
    assign n1169 = n759 ? n329 : m_a1[27];   // insn_decoder.v(198)
    assign n1171 = n759 ? n330 : m_a1[26];   // insn_decoder.v(198)
    assign n1173 = n759 ? n331 : m_a1[25];   // insn_decoder.v(198)
    assign n1175 = n759 ? n332 : m_a1[24];   // insn_decoder.v(198)
    assign n1177 = n759 ? n333 : m_a1[23];   // insn_decoder.v(198)
    assign n1179 = n759 ? n334 : m_a1[22];   // insn_decoder.v(198)
    assign n1181 = n759 ? n335 : m_a1[21];   // insn_decoder.v(198)
    assign n1183 = n759 ? n336 : m_a1[20];   // insn_decoder.v(198)
    assign n1185 = n759 ? n337 : m_a1[19];   // insn_decoder.v(198)
    assign n1187 = n759 ? n338 : m_a1[18];   // insn_decoder.v(198)
    assign n1189 = n759 ? n339 : m_a1[17];   // insn_decoder.v(198)
    assign n1191 = n759 ? n340 : m_a1[16];   // insn_decoder.v(198)
    assign n1193 = n759 ? n341 : m_a1[15];   // insn_decoder.v(198)
    assign n1195 = n759 ? n342 : m_a1[14];   // insn_decoder.v(198)
    assign n1197 = n759 ? n343 : m_a1[13];   // insn_decoder.v(198)
    assign n1199 = n759 ? n344 : m_a1[12];   // insn_decoder.v(198)
    assign n1201 = n759 ? n345 : m_a1[11];   // insn_decoder.v(198)
    assign n1203 = n759 ? n346 : m_a1[10];   // insn_decoder.v(198)
    assign n1205 = n759 ? n347 : m_a1[9];   // insn_decoder.v(198)
    assign n1207 = n759 ? n348 : m_a1[8];   // insn_decoder.v(198)
    assign n1209 = n759 ? n349 : m_a1[7];   // insn_decoder.v(198)
    assign n1211 = n759 ? n350 : m_a1[6];   // insn_decoder.v(198)
    assign n1213 = n759 ? n351 : m_a1[5];   // insn_decoder.v(198)
    assign n1215 = n759 ? n352 : m_a1[4];   // insn_decoder.v(198)
    assign n1217 = n759 ? n353 : m_a1[3];   // insn_decoder.v(198)
    assign n1219 = n759 ? n354 : m_a1[2];   // insn_decoder.v(198)
    assign n1221 = n759 ? n355 : m_a1[1];   // insn_decoder.v(198)
    assign n1223 = n759 ? n356 : m_a1[0];   // insn_decoder.v(198)
    or (n1224, n524, n657, n660, n663, n666, n669, n672, n675, 
        n678, n681, n684, n687, n690, n693, n696, n699, n702, 
        n705, n708, n711, n714, n717, n720, n723, n726, n729, 
        n732, n735, n738, n741, n744, n747, n750, n753, n756, 
        n765, n768, n770) ;   // insn_decoder.v(198)
    Select_3 Select_1220 (.sel({n1224, n759, n762}), .data({m_a2[31], 
            n357, n460}), .o(n1225));   // insn_decoder.v(198)
    Select_3 Select_1222 (.sel({n1224, n759, n762}), .data({m_a2[30], 
            n358, n461}), .o(n1227));   // insn_decoder.v(198)
    Select_3 Select_1224 (.sel({n1224, n759, n762}), .data({m_a2[29], 
            n359, n462}), .o(n1229));   // insn_decoder.v(198)
    Select_3 Select_1226 (.sel({n1224, n759, n762}), .data({m_a2[28], 
            n360, n463}), .o(n1231));   // insn_decoder.v(198)
    Select_3 Select_1228 (.sel({n1224, n759, n762}), .data({m_a2[27], 
            n361, n464}), .o(n1233));   // insn_decoder.v(198)
    Select_3 Select_1230 (.sel({n1224, n759, n762}), .data({m_a2[26], 
            n362, n465}), .o(n1235));   // insn_decoder.v(198)
    Select_3 Select_1232 (.sel({n1224, n759, n762}), .data({m_a2[25], 
            n363, n466}), .o(n1237));   // insn_decoder.v(198)
    Select_3 Select_1234 (.sel({n1224, n759, n762}), .data({m_a2[24], 
            n364, n467}), .o(n1239));   // insn_decoder.v(198)
    Select_3 Select_1236 (.sel({n1224, n759, n762}), .data({m_a2[23], 
            n365, n468}), .o(n1241));   // insn_decoder.v(198)
    Select_3 Select_1238 (.sel({n1224, n759, n762}), .data({m_a2[22], 
            n366, n469}), .o(n1243));   // insn_decoder.v(198)
    Select_3 Select_1240 (.sel({n1224, n759, n762}), .data({m_a2[21], 
            n367, n470}), .o(n1245));   // insn_decoder.v(198)
    Select_3 Select_1242 (.sel({n1224, n759, n762}), .data({m_a2[20], 
            n368, n471}), .o(n1247));   // insn_decoder.v(198)
    Select_3 Select_1244 (.sel({n1224, n759, n762}), .data({m_a2[19], 
            n369, n472}), .o(n1249));   // insn_decoder.v(198)
    Select_3 Select_1246 (.sel({n1224, n759, n762}), .data({m_a2[18], 
            n370, n473}), .o(n1251));   // insn_decoder.v(198)
    Select_3 Select_1248 (.sel({n1224, n759, n762}), .data({m_a2[17], 
            n371, n474}), .o(n1253));   // insn_decoder.v(198)
    Select_3 Select_1250 (.sel({n1224, n759, n762}), .data({m_a2[16], 
            n372, n475}), .o(n1255));   // insn_decoder.v(198)
    Select_3 Select_1252 (.sel({n1224, n759, n762}), .data({m_a2[15], 
            n373, n476}), .o(n1257));   // insn_decoder.v(198)
    Select_3 Select_1254 (.sel({n1224, n759, n762}), .data({m_a2[14], 
            n374, n477}), .o(n1259));   // insn_decoder.v(198)
    Select_3 Select_1256 (.sel({n1224, n759, n762}), .data({m_a2[13], 
            n375, n478}), .o(n1261));   // insn_decoder.v(198)
    Select_3 Select_1258 (.sel({n1224, n759, n762}), .data({m_a2[12], 
            n376, n479}), .o(n1263));   // insn_decoder.v(198)
    Select_3 Select_1260 (.sel({n1224, n759, n762}), .data({m_a2[11], 
            n377, n480}), .o(n1265));   // insn_decoder.v(198)
    Select_3 Select_1262 (.sel({n1224, n759, n762}), .data({m_a2[10], 
            n378, n481}), .o(n1267));   // insn_decoder.v(198)
    Select_3 Select_1264 (.sel({n1224, n759, n762}), .data({m_a2[9], 
            n379, n482}), .o(n1269));   // insn_decoder.v(198)
    Select_3 Select_1266 (.sel({n1224, n759, n762}), .data({m_a2[8], 
            n380, n483}), .o(n1271));   // insn_decoder.v(198)
    Select_3 Select_1268 (.sel({n1224, n759, n762}), .data({m_a2[7], 
            n381, n484}), .o(n1273));   // insn_decoder.v(198)
    Select_3 Select_1270 (.sel({n1224, n759, n762}), .data({m_a2[6], 
            n382, n485}), .o(n1275));   // insn_decoder.v(198)
    Select_3 Select_1272 (.sel({n1224, n759, n762}), .data({m_a2[5], 
            n383, n486}), .o(n1277));   // insn_decoder.v(198)
    Select_3 Select_1274 (.sel({n1224, n759, n762}), .data({m_a2[4], 
            n384, n487}), .o(n1279));   // insn_decoder.v(198)
    Select_3 Select_1276 (.sel({n1224, n759, n762}), .data({m_a2[3], 
            n385, n488}), .o(n1281));   // insn_decoder.v(198)
    Select_3 Select_1278 (.sel({n1224, n759, n762}), .data({m_a2[2], 
            n386, n489}), .o(n1283));   // insn_decoder.v(198)
    Select_3 Select_1280 (.sel({n1224, n759, n762}), .data({m_a2[1], 
            n387, n490}), .o(n1285));   // insn_decoder.v(198)
    Select_3 Select_1282 (.sel({n1224, n759, n762}), .data({m_a2[0], 
            n388, n491}), .o(n1287));   // insn_decoder.v(198)
    or (n1288, n524, n657, n660, n663, n666, n669, n672, n675, 
            n678, n681, n684, n687, n690, n693, n696, n699, 
            n702, n705, n708, n711, n714, n717, n720, n723, 
            n726, n729, n732, n735, n738, n741, n744, n747, 
            n750, n753, n756, n759, n762, n770) ;   // insn_decoder.v(198)
    Select_3 Select_1284 (.sel({n1288, n765, n768}), .data({n48, 1'b0, 
            n513}), .o(n1289));   // insn_decoder.v(198)
    assign n1291 = n768 ? n514 : n49;   // insn_decoder.v(198)
    assign n1292 = set_delay ? 1'b0 : n1056;   // insn_decoder.v(555)
    assign n1293 = set_delay ? 1'b0 : n1059;   // insn_decoder.v(555)
    assign n1294 = set_delay ? 1'b1 : n1062;   // insn_decoder.v(555)
    assign n1295 = set_delay ? 1'b0 : n1065;   // insn_decoder.v(555)
    assign n1296 = set_delay ? 1'b0 : n1068;   // insn_decoder.v(555)
    assign n1297 = set_delay ? 1'b0 : n1071;   // insn_decoder.v(555)
    assign n1298 = set_delay ? 1'b0 : n1074;   // insn_decoder.v(555)
    assign n1299 = set_delay ? 1'b0 : n1077;   // insn_decoder.v(555)
    assign n1300 = set_delay ? 1'b1 : n1080;   // insn_decoder.v(555)
    assign n1301 = set_delay ? 1'b0 : n1083;   // insn_decoder.v(555)
    assign n1302 = set_delay ? 1'b0 : set_delay;   // insn_decoder.v(555)
    or (n1304, n59, imm_action[1], imm_action[0]) ;   // insn_decoder.v(561)
    or (n1305, imm_action[2], imm_action[1], imm_action[0]) ;   // insn_decoder.v(561)
    and (n1306, n1304, n1305) ;   // insn_decoder.v(561)
    or (n1308, n644, state1[6], state1[5], state1[4], state1[3], 
        state1[2], state1[1], state1[0]) ;   // insn_decoder.v(562)
    or (n1311, n644, state1[6], state1[5], state1[4], state1[3], 
        state1[2], state1[1], n525) ;   // insn_decoder.v(562)
    and (n1312, n1308, n1311) ;   // insn_decoder.v(562)
    assign n1313 = imm_action[1] ? 1'b0 : n872;   // insn_decoder.v(563)
    assign n1314 = imm_action[0] ? 1'b0 : n869;   // insn_decoder.v(566)
    or (n1324, n391, n395) ;   // insn_decoder.v(580)
    assign n1325 = n1324 ? 1'b0 : old_pass_imm;   // insn_decoder.v(587)
    assign n1326 = n1324 ? 1'b0 : old_fetch_imm;   // insn_decoder.v(587)
    not (n1327, n1324) ;   // insn_decoder.v(587)
    assign n1328 = n1324 ? 1'b1 : old_pcincr_imm;   // insn_decoder.v(587)
    assign n1329 = n1324 ? 1'b1 : old_state1_imm[7];   // insn_decoder.v(587)
    assign n1330 = n1324 ? 1'b0 : old_state1_imm[6];   // insn_decoder.v(587)
    assign n1331 = n1324 ? 1'b0 : old_state1_imm[5];   // insn_decoder.v(587)
    assign n1332 = n1324 ? 1'b0 : old_state1_imm[4];   // insn_decoder.v(587)
    assign n1333 = n1324 ? 1'b0 : old_state1_imm[3];   // insn_decoder.v(587)
    assign n1334 = n1324 ? 1'b0 : old_state1_imm[2];   // insn_decoder.v(587)
    assign n1335 = n1324 ? 1'b0 : old_state1_imm[1];   // insn_decoder.v(587)
    assign n1336 = n1324 ? 1'b1 : old_state1_imm[0];   // insn_decoder.v(587)
    assign n1337 = n1324 ? n936 : 1'b0;   // insn_decoder.v(587)
    assign n1338 = n1324 ? n939 : 1'b0;   // insn_decoder.v(587)
    assign n1339 = n1324 ? n942 : 1'b0;   // insn_decoder.v(587)
    assign n1343 = n1342 ? old_state1_imm[7] : n1294;   // insn_decoder.v(596)
    assign n1344 = n1342 ? old_state1_imm[6] : n1295;   // insn_decoder.v(596)
    assign n1345 = n1342 ? old_state1_imm[5] : n1296;   // insn_decoder.v(596)
    assign n1346 = n1342 ? old_state1_imm[4] : n1297;   // insn_decoder.v(596)
    assign n1347 = n1342 ? old_state1_imm[3] : n1298;   // insn_decoder.v(596)
    assign n1348 = n1342 ? old_state1_imm[2] : n1299;   // insn_decoder.v(596)
    assign n1349 = n1342 ? old_state1_imm[1] : n1300;   // insn_decoder.v(596)
    assign n1350 = n1342 ? old_state1_imm[0] : n1301;   // insn_decoder.v(596)
    assign n1351 = n1342 ? old_pass_imm : n1289;   // insn_decoder.v(596)
    assign n1352 = n1342 ? old_fetch_imm : n1292;   // insn_decoder.v(596)
    assign n1353 = n1342 ? old_pcincr_imm : n1293;   // insn_decoder.v(596)
    assign n1354 = n1342 ? 1'b1 : n1291;   // insn_decoder.v(596)
    assign n1355 = n1342 ? 1'b0 : n936;   // insn_decoder.v(596)
    assign n1356 = n1342 ? 1'b0 : n939;   // insn_decoder.v(596)
    assign n1357 = n1342 ? 1'b0 : n942;   // insn_decoder.v(596)
    assign n1358 = n1316 ? n1325 : n1351;   // insn_decoder.v(596)
    assign n1359 = n1316 ? n1326 : n1352;   // insn_decoder.v(596)
    assign n1360 = n1316 ? n1327 : n1354;   // insn_decoder.v(596)
    assign n1361 = n1316 ? n1328 : n1353;   // insn_decoder.v(596)
    assign n1362 = n1316 ? n1329 : n1343;   // insn_decoder.v(596)
    assign n1363 = n1316 ? n1330 : n1344;   // insn_decoder.v(596)
    assign n1364 = n1316 ? n1331 : n1345;   // insn_decoder.v(596)
    assign n1365 = n1316 ? n1332 : n1346;   // insn_decoder.v(596)
    assign n1366 = n1316 ? n1333 : n1347;   // insn_decoder.v(596)
    assign n1367 = n1316 ? n1334 : n1348;   // insn_decoder.v(596)
    assign n1368 = n1316 ? n1335 : n1349;   // insn_decoder.v(596)
    assign n1369 = n1316 ? n1336 : n1350;   // insn_decoder.v(596)
    assign n1370 = n1316 ? n1337 : n1355;   // insn_decoder.v(596)
    assign n1371 = n1316 ? n1338 : n1356;   // insn_decoder.v(596)
    assign n1372 = n1316 ? n1339 : n1357;   // insn_decoder.v(596)
    assign n1373 = n1312 ? n1314 : n869;   // insn_decoder.v(579)
    assign n1374 = n1312 ? n1313 : n872;   // insn_decoder.v(579)
    assign n1375 = n1312 ? state1[7] : old_state1_imm[7];   // insn_decoder.v(579)
    assign n1376 = n1312 ? state1[6] : old_state1_imm[6];   // insn_decoder.v(579)
    assign n1377 = n1312 ? state1[5] : old_state1_imm[5];   // insn_decoder.v(579)
    assign n1378 = n1312 ? state1[4] : old_state1_imm[4];   // insn_decoder.v(579)
    assign n1379 = n1312 ? state1[3] : old_state1_imm[3];   // insn_decoder.v(579)
    assign n1380 = n1312 ? state1[2] : old_state1_imm[2];   // insn_decoder.v(579)
    assign n1381 = n1312 ? state1[1] : old_state1_imm[1];   // insn_decoder.v(579)
    assign n1382 = n1312 ? state1[0] : old_state1_imm[0];   // insn_decoder.v(579)
    assign n1383 = n1312 ? d_pass : old_pass_imm;   // insn_decoder.v(579)
    assign n1384 = n1312 ? fetch : old_fetch_imm;   // insn_decoder.v(579)
    assign n1385 = n1312 ? d_pcincr : old_pcincr_imm;   // insn_decoder.v(579)
    assign n1386 = n1312 ? 1'b0 : n1358;   // insn_decoder.v(579)
    assign n1387 = n1312 ? 1'b0 : n1359;   // insn_decoder.v(579)
    assign n1388 = n1312 ? 1'b0 : n1360;   // insn_decoder.v(579)
    assign n1389 = n1312 ? 1'b1 : n1361;   // insn_decoder.v(579)
    assign n1390 = n1312 ? 1'b1 : n1362;   // insn_decoder.v(579)
    assign n1391 = n1312 ? 1'b0 : n1363;   // insn_decoder.v(579)
    assign n1392 = n1312 ? 1'b0 : n1364;   // insn_decoder.v(579)
    assign n1393 = n1312 ? 1'b0 : n1365;   // insn_decoder.v(579)
    assign n1394 = n1312 ? 1'b0 : n1366;   // insn_decoder.v(579)
    assign n1395 = n1312 ? 1'b0 : n1367;   // insn_decoder.v(579)
    assign n1396 = n1312 ? 1'b0 : n1368;   // insn_decoder.v(579)
    assign n1397 = n1312 ? 1'b0 : n1369;   // insn_decoder.v(579)
    assign n1398 = n1312 ? n936 : n1370;   // insn_decoder.v(579)
    assign n1399 = n1312 ? n939 : n1371;   // insn_decoder.v(579)
    assign n1400 = n1312 ? n942 : n1372;   // insn_decoder.v(579)
    assign n1401 = n1306 ? n1373 : n869;   // insn_decoder.v(561)
    assign n1402 = n1306 ? n1374 : n872;   // insn_decoder.v(561)
    assign n1403 = n1306 ? n1375 : old_state1_imm[7];   // insn_decoder.v(561)
    assign n1404 = n1306 ? n1376 : old_state1_imm[6];   // insn_decoder.v(561)
    assign n1405 = n1306 ? n1377 : old_state1_imm[5];   // insn_decoder.v(561)
    assign n1406 = n1306 ? n1378 : old_state1_imm[4];   // insn_decoder.v(561)
    assign n1407 = n1306 ? n1379 : old_state1_imm[3];   // insn_decoder.v(561)
    assign n1408 = n1306 ? n1380 : old_state1_imm[2];   // insn_decoder.v(561)
    assign n1409 = n1306 ? n1381 : old_state1_imm[1];   // insn_decoder.v(561)
    assign n1410 = n1306 ? n1382 : old_state1_imm[0];   // insn_decoder.v(561)
    assign n1411 = n1306 ? n1383 : old_pass_imm;   // insn_decoder.v(561)
    assign n1412 = n1306 ? n1384 : old_fetch_imm;   // insn_decoder.v(561)
    assign n1413 = n1306 ? n1385 : old_pcincr_imm;   // insn_decoder.v(561)
    assign n1414 = n1306 ? n1386 : n1289;   // insn_decoder.v(561)
    assign n1415 = n1306 ? n1387 : n1292;   // insn_decoder.v(561)
    assign n1416 = n1306 ? n1388 : n1291;   // insn_decoder.v(561)
    assign n1417 = n1306 ? n1389 : n1293;   // insn_decoder.v(561)
    assign n1418 = n1306 ? n1390 : n1294;   // insn_decoder.v(561)
    assign n1419 = n1306 ? n1391 : n1295;   // insn_decoder.v(561)
    assign n1420 = n1306 ? n1392 : n1296;   // insn_decoder.v(561)
    assign n1421 = n1306 ? n1393 : n1297;   // insn_decoder.v(561)
    assign n1422 = n1306 ? n1394 : n1298;   // insn_decoder.v(561)
    assign n1423 = n1306 ? n1395 : n1299;   // insn_decoder.v(561)
    assign n1424 = n1306 ? n1396 : n1300;   // insn_decoder.v(561)
    assign n1425 = n1306 ? n1397 : n1301;   // insn_decoder.v(561)
    assign n1426 = n1306 ? n1398 : n936;   // insn_decoder.v(561)
    assign n1427 = n1306 ? n1399 : n939;   // insn_decoder.v(561)
    assign n1428 = n1306 ? n1400 : n942;   // insn_decoder.v(561)
    and (n1429, hazard, reg_fetch) ;   // insn_decoder.v(606)
    assign n1430 = n1429 ? d_pcincr : old_pcincr_hz;   // insn_decoder.v(606)
    assign n1431 = n1429 ? d_pass : old_pass_hz;   // insn_decoder.v(606)
    assign n1432 = n1429 ? fetch : old_fetch_hz;   // insn_decoder.v(606)
    assign n1433 = n1429 ? state1[7] : old_state1_hz[7];   // insn_decoder.v(606)
    assign n1434 = n1429 ? state1[6] : old_state1_hz[6];   // insn_decoder.v(606)
    assign n1435 = n1429 ? state1[5] : old_state1_hz[5];   // insn_decoder.v(606)
    assign n1436 = n1429 ? state1[4] : old_state1_hz[4];   // insn_decoder.v(606)
    assign n1437 = n1429 ? state1[3] : old_state1_hz[3];   // insn_decoder.v(606)
    assign n1438 = n1429 ? state1[2] : old_state1_hz[2];   // insn_decoder.v(606)
    assign n1439 = n1429 ? state1[1] : old_state1_hz[1];   // insn_decoder.v(606)
    assign n1440 = n1429 ? state1[0] : old_state1_hz[0];   // insn_decoder.v(606)
    assign n1441 = n1429 ? 1'b0 : n1417;   // insn_decoder.v(606)
    assign n1442 = n1429 ? 1'b0 : n1414;   // insn_decoder.v(606)
    assign n1443 = n1429 ? 1'b0 : n1415;   // insn_decoder.v(606)
    assign n1444 = n1429 ? 1'b0 : n1416;   // insn_decoder.v(606)
    assign n1445 = n1429 ? 1'b1 : n1418;   // insn_decoder.v(606)
    assign n1446 = n1429 ? 1'b0 : n1419;   // insn_decoder.v(606)
    assign n1447 = n1429 ? 1'b0 : n1420;   // insn_decoder.v(606)
    assign n1448 = n1429 ? 1'b0 : n1421;   // insn_decoder.v(606)
    assign n1449 = n1429 ? 1'b0 : n1422;   // insn_decoder.v(606)
    assign n1450 = n1429 ? 1'b0 : n1423;   // insn_decoder.v(606)
    assign n1451 = n1429 ? 1'b1 : n1424;   // insn_decoder.v(606)
    assign n1452 = n1429 ? 1'b1 : n1425;   // insn_decoder.v(606)
    assign n1453 = r_to_mem[0] ? r1[31] : n1161;   // insn_decoder.v(621)
    assign n1454 = r_to_mem[0] ? r1[30] : n1163;   // insn_decoder.v(621)
    assign n1455 = r_to_mem[0] ? r1[29] : n1165;   // insn_decoder.v(621)
    assign n1456 = r_to_mem[0] ? r1[28] : n1167;   // insn_decoder.v(621)
    assign n1457 = r_to_mem[0] ? r1[27] : n1169;   // insn_decoder.v(621)
    assign n1458 = r_to_mem[0] ? r1[26] : n1171;   // insn_decoder.v(621)
    assign n1459 = r_to_mem[0] ? r1[25] : n1173;   // insn_decoder.v(621)
    assign n1460 = r_to_mem[0] ? r1[24] : n1175;   // insn_decoder.v(621)
    assign n1461 = r_to_mem[0] ? r1[23] : n1177;   // insn_decoder.v(621)
    assign n1462 = r_to_mem[0] ? r1[22] : n1179;   // insn_decoder.v(621)
    assign n1463 = r_to_mem[0] ? r1[21] : n1181;   // insn_decoder.v(621)
    assign n1464 = r_to_mem[0] ? r1[20] : n1183;   // insn_decoder.v(621)
    assign n1465 = r_to_mem[0] ? r1[19] : n1185;   // insn_decoder.v(621)
    assign n1466 = r_to_mem[0] ? r1[18] : n1187;   // insn_decoder.v(621)
    assign n1467 = r_to_mem[0] ? r1[17] : n1189;   // insn_decoder.v(621)
    assign n1468 = r_to_mem[0] ? r1[16] : n1191;   // insn_decoder.v(621)
    assign n1469 = r_to_mem[0] ? r1[15] : n1193;   // insn_decoder.v(621)
    assign n1470 = r_to_mem[0] ? r1[14] : n1195;   // insn_decoder.v(621)
    assign n1471 = r_to_mem[0] ? r1[13] : n1197;   // insn_decoder.v(621)
    assign n1472 = r_to_mem[0] ? r1[12] : n1199;   // insn_decoder.v(621)
    assign n1473 = r_to_mem[0] ? r1[11] : n1201;   // insn_decoder.v(621)
    assign n1474 = r_to_mem[0] ? r1[10] : n1203;   // insn_decoder.v(621)
    assign n1475 = r_to_mem[0] ? r1[9] : n1205;   // insn_decoder.v(621)
    assign n1476 = r_to_mem[0] ? r1[8] : n1207;   // insn_decoder.v(621)
    assign n1477 = r_to_mem[0] ? r1[7] : n1209;   // insn_decoder.v(621)
    assign n1478 = r_to_mem[0] ? r1[6] : n1211;   // insn_decoder.v(621)
    assign n1479 = r_to_mem[0] ? r1[5] : n1213;   // insn_decoder.v(621)
    assign n1480 = r_to_mem[0] ? r1[4] : n1215;   // insn_decoder.v(621)
    assign n1481 = r_to_mem[0] ? r1[3] : n1217;   // insn_decoder.v(621)
    assign n1482 = r_to_mem[0] ? r1[2] : n1219;   // insn_decoder.v(621)
    assign n1483 = r_to_mem[0] ? r1[1] : n1221;   // insn_decoder.v(621)
    assign n1484 = r_to_mem[0] ? r1[0] : n1223;   // insn_decoder.v(621)
    assign n1485 = r_to_mem[0] ? n1097 : r1[31];   // insn_decoder.v(621)
    assign n1486 = r_to_mem[0] ? n1099 : r1[30];   // insn_decoder.v(621)
    assign n1487 = r_to_mem[0] ? n1101 : r1[29];   // insn_decoder.v(621)
    assign n1488 = r_to_mem[0] ? n1103 : r1[28];   // insn_decoder.v(621)
    assign n1489 = r_to_mem[0] ? n1105 : r1[27];   // insn_decoder.v(621)
    assign n1490 = r_to_mem[0] ? n1107 : r1[26];   // insn_decoder.v(621)
    assign n1491 = r_to_mem[0] ? n1109 : r1[25];   // insn_decoder.v(621)
    assign n1492 = r_to_mem[0] ? n1111 : r1[24];   // insn_decoder.v(621)
    assign n1493 = r_to_mem[0] ? n1113 : r1[23];   // insn_decoder.v(621)
    assign n1494 = r_to_mem[0] ? n1115 : r1[22];   // insn_decoder.v(621)
    assign n1495 = r_to_mem[0] ? n1117 : r1[21];   // insn_decoder.v(621)
    assign n1496 = r_to_mem[0] ? n1119 : r1[20];   // insn_decoder.v(621)
    assign n1497 = r_to_mem[0] ? n1121 : r1[19];   // insn_decoder.v(621)
    assign n1498 = r_to_mem[0] ? n1123 : r1[18];   // insn_decoder.v(621)
    assign n1499 = r_to_mem[0] ? n1125 : r1[17];   // insn_decoder.v(621)
    assign n1500 = r_to_mem[0] ? n1127 : r1[16];   // insn_decoder.v(621)
    assign n1501 = r_to_mem[0] ? n1129 : r1[15];   // insn_decoder.v(621)
    assign n1502 = r_to_mem[0] ? n1131 : r1[14];   // insn_decoder.v(621)
    assign n1503 = r_to_mem[0] ? n1133 : r1[13];   // insn_decoder.v(621)
    assign n1504 = r_to_mem[0] ? n1135 : r1[12];   // insn_decoder.v(621)
    assign n1505 = r_to_mem[0] ? n1137 : r1[11];   // insn_decoder.v(621)
    assign n1506 = r_to_mem[0] ? n1139 : r1[10];   // insn_decoder.v(621)
    assign n1507 = r_to_mem[0] ? n1141 : r1[9];   // insn_decoder.v(621)
    assign n1508 = r_to_mem[0] ? n1143 : r1[8];   // insn_decoder.v(621)
    assign n1509 = r_to_mem[0] ? n1145 : r1[7];   // insn_decoder.v(621)
    assign n1510 = r_to_mem[0] ? n1147 : r1[6];   // insn_decoder.v(621)
    assign n1511 = r_to_mem[0] ? n1149 : r1[5];   // insn_decoder.v(621)
    assign n1512 = r_to_mem[0] ? n1151 : r1[4];   // insn_decoder.v(621)
    assign n1513 = r_to_mem[0] ? n1153 : r1[3];   // insn_decoder.v(621)
    assign n1514 = r_to_mem[0] ? n1155 : r1[2];   // insn_decoder.v(621)
    assign n1515 = r_to_mem[0] ? n1157 : r1[1];   // insn_decoder.v(621)
    assign n1516 = r_to_mem[0] ? n1159 : r1[0];   // insn_decoder.v(621)
    assign n1517 = r_read[0] ? n1453 : n1161;   // insn_decoder.v(619)
    assign n1518 = r_read[0] ? n1454 : n1163;   // insn_decoder.v(619)
    assign n1519 = r_read[0] ? n1455 : n1165;   // insn_decoder.v(619)
    assign n1520 = r_read[0] ? n1456 : n1167;   // insn_decoder.v(619)
    assign n1521 = r_read[0] ? n1457 : n1169;   // insn_decoder.v(619)
    assign n1522 = r_read[0] ? n1458 : n1171;   // insn_decoder.v(619)
    assign n1523 = r_read[0] ? n1459 : n1173;   // insn_decoder.v(619)
    assign n1524 = r_read[0] ? n1460 : n1175;   // insn_decoder.v(619)
    assign n1525 = r_read[0] ? n1461 : n1177;   // insn_decoder.v(619)
    assign n1526 = r_read[0] ? n1462 : n1179;   // insn_decoder.v(619)
    assign n1527 = r_read[0] ? n1463 : n1181;   // insn_decoder.v(619)
    assign n1528 = r_read[0] ? n1464 : n1183;   // insn_decoder.v(619)
    assign n1529 = r_read[0] ? n1465 : n1185;   // insn_decoder.v(619)
    assign n1530 = r_read[0] ? n1466 : n1187;   // insn_decoder.v(619)
    assign n1531 = r_read[0] ? n1467 : n1189;   // insn_decoder.v(619)
    assign n1532 = r_read[0] ? n1468 : n1191;   // insn_decoder.v(619)
    assign n1533 = r_read[0] ? n1469 : n1193;   // insn_decoder.v(619)
    assign n1534 = r_read[0] ? n1470 : n1195;   // insn_decoder.v(619)
    assign n1535 = r_read[0] ? n1471 : n1197;   // insn_decoder.v(619)
    assign n1536 = r_read[0] ? n1472 : n1199;   // insn_decoder.v(619)
    assign n1537 = r_read[0] ? n1473 : n1201;   // insn_decoder.v(619)
    assign n1538 = r_read[0] ? n1474 : n1203;   // insn_decoder.v(619)
    assign n1539 = r_read[0] ? n1475 : n1205;   // insn_decoder.v(619)
    assign n1540 = r_read[0] ? n1476 : n1207;   // insn_decoder.v(619)
    assign n1541 = r_read[0] ? n1477 : n1209;   // insn_decoder.v(619)
    assign n1542 = r_read[0] ? n1478 : n1211;   // insn_decoder.v(619)
    assign n1543 = r_read[0] ? n1479 : n1213;   // insn_decoder.v(619)
    assign n1544 = r_read[0] ? n1480 : n1215;   // insn_decoder.v(619)
    assign n1545 = r_read[0] ? n1481 : n1217;   // insn_decoder.v(619)
    assign n1546 = r_read[0] ? n1482 : n1219;   // insn_decoder.v(619)
    assign n1547 = r_read[0] ? n1483 : n1221;   // insn_decoder.v(619)
    assign n1548 = r_read[0] ? n1484 : n1223;   // insn_decoder.v(619)
    assign n1549 = r_read[0] ? n1485 : n1097;   // insn_decoder.v(619)
    assign n1550 = r_read[0] ? n1486 : n1099;   // insn_decoder.v(619)
    assign n1551 = r_read[0] ? n1487 : n1101;   // insn_decoder.v(619)
    assign n1552 = r_read[0] ? n1488 : n1103;   // insn_decoder.v(619)
    assign n1553 = r_read[0] ? n1489 : n1105;   // insn_decoder.v(619)
    assign n1554 = r_read[0] ? n1490 : n1107;   // insn_decoder.v(619)
    assign n1555 = r_read[0] ? n1491 : n1109;   // insn_decoder.v(619)
    assign n1556 = r_read[0] ? n1492 : n1111;   // insn_decoder.v(619)
    assign n1557 = r_read[0] ? n1493 : n1113;   // insn_decoder.v(619)
    assign n1558 = r_read[0] ? n1494 : n1115;   // insn_decoder.v(619)
    assign n1559 = r_read[0] ? n1495 : n1117;   // insn_decoder.v(619)
    assign n1560 = r_read[0] ? n1496 : n1119;   // insn_decoder.v(619)
    assign n1561 = r_read[0] ? n1497 : n1121;   // insn_decoder.v(619)
    assign n1562 = r_read[0] ? n1498 : n1123;   // insn_decoder.v(619)
    assign n1563 = r_read[0] ? n1499 : n1125;   // insn_decoder.v(619)
    assign n1564 = r_read[0] ? n1500 : n1127;   // insn_decoder.v(619)
    assign n1565 = r_read[0] ? n1501 : n1129;   // insn_decoder.v(619)
    assign n1566 = r_read[0] ? n1502 : n1131;   // insn_decoder.v(619)
    assign n1567 = r_read[0] ? n1503 : n1133;   // insn_decoder.v(619)
    assign n1568 = r_read[0] ? n1504 : n1135;   // insn_decoder.v(619)
    assign n1569 = r_read[0] ? n1505 : n1137;   // insn_decoder.v(619)
    assign n1570 = r_read[0] ? n1506 : n1139;   // insn_decoder.v(619)
    assign n1571 = r_read[0] ? n1507 : n1141;   // insn_decoder.v(619)
    assign n1572 = r_read[0] ? n1508 : n1143;   // insn_decoder.v(619)
    assign n1573 = r_read[0] ? n1509 : n1145;   // insn_decoder.v(619)
    assign n1574 = r_read[0] ? n1510 : n1147;   // insn_decoder.v(619)
    assign n1575 = r_read[0] ? n1511 : n1149;   // insn_decoder.v(619)
    assign n1576 = r_read[0] ? n1512 : n1151;   // insn_decoder.v(619)
    assign n1577 = r_read[0] ? n1513 : n1153;   // insn_decoder.v(619)
    assign n1578 = r_read[0] ? n1514 : n1155;   // insn_decoder.v(619)
    assign n1579 = r_read[0] ? n1515 : n1157;   // insn_decoder.v(619)
    assign n1580 = r_read[0] ? n1516 : n1159;   // insn_decoder.v(619)
    assign n1581 = r_to_mem[1] ? r2[31] : n1225;   // insn_decoder.v(625)
    assign n1582 = r_to_mem[1] ? r2[30] : n1227;   // insn_decoder.v(625)
    assign n1583 = r_to_mem[1] ? r2[29] : n1229;   // insn_decoder.v(625)
    assign n1584 = r_to_mem[1] ? r2[28] : n1231;   // insn_decoder.v(625)
    assign n1585 = r_to_mem[1] ? r2[27] : n1233;   // insn_decoder.v(625)
    assign n1586 = r_to_mem[1] ? r2[26] : n1235;   // insn_decoder.v(625)
    assign n1587 = r_to_mem[1] ? r2[25] : n1237;   // insn_decoder.v(625)
    assign n1588 = r_to_mem[1] ? r2[24] : n1239;   // insn_decoder.v(625)
    assign n1589 = r_to_mem[1] ? r2[23] : n1241;   // insn_decoder.v(625)
    assign n1590 = r_to_mem[1] ? r2[22] : n1243;   // insn_decoder.v(625)
    assign n1591 = r_to_mem[1] ? r2[21] : n1245;   // insn_decoder.v(625)
    assign n1592 = r_to_mem[1] ? r2[20] : n1247;   // insn_decoder.v(625)
    assign n1593 = r_to_mem[1] ? r2[19] : n1249;   // insn_decoder.v(625)
    assign n1594 = r_to_mem[1] ? r2[18] : n1251;   // insn_decoder.v(625)
    assign n1595 = r_to_mem[1] ? r2[17] : n1253;   // insn_decoder.v(625)
    assign n1596 = r_to_mem[1] ? r2[16] : n1255;   // insn_decoder.v(625)
    assign n1597 = r_to_mem[1] ? r2[15] : n1257;   // insn_decoder.v(625)
    assign n1598 = r_to_mem[1] ? r2[14] : n1259;   // insn_decoder.v(625)
    assign n1599 = r_to_mem[1] ? r2[13] : n1261;   // insn_decoder.v(625)
    assign n1600 = r_to_mem[1] ? r2[12] : n1263;   // insn_decoder.v(625)
    assign n1601 = r_to_mem[1] ? r2[11] : n1265;   // insn_decoder.v(625)
    assign n1602 = r_to_mem[1] ? r2[10] : n1267;   // insn_decoder.v(625)
    assign n1603 = r_to_mem[1] ? r2[9] : n1269;   // insn_decoder.v(625)
    assign n1604 = r_to_mem[1] ? r2[8] : n1271;   // insn_decoder.v(625)
    assign n1605 = r_to_mem[1] ? r2[7] : n1273;   // insn_decoder.v(625)
    assign n1606 = r_to_mem[1] ? r2[6] : n1275;   // insn_decoder.v(625)
    assign n1607 = r_to_mem[1] ? r2[5] : n1277;   // insn_decoder.v(625)
    assign n1608 = r_to_mem[1] ? r2[4] : n1279;   // insn_decoder.v(625)
    assign n1609 = r_to_mem[1] ? r2[3] : n1281;   // insn_decoder.v(625)
    assign n1610 = r_to_mem[1] ? r2[2] : n1283;   // insn_decoder.v(625)
    assign n1611 = r_to_mem[1] ? r2[1] : n1285;   // insn_decoder.v(625)
    assign n1612 = r_to_mem[1] ? r2[0] : n1287;   // insn_decoder.v(625)
    assign n1613 = r_to_mem[1] ? n960 : r2[31];   // insn_decoder.v(625)
    assign n1614 = r_to_mem[1] ? n963 : r2[30];   // insn_decoder.v(625)
    assign n1615 = r_to_mem[1] ? n966 : r2[29];   // insn_decoder.v(625)
    assign n1616 = r_to_mem[1] ? n969 : r2[28];   // insn_decoder.v(625)
    assign n1617 = r_to_mem[1] ? n972 : r2[27];   // insn_decoder.v(625)
    assign n1618 = r_to_mem[1] ? n975 : r2[26];   // insn_decoder.v(625)
    assign n1619 = r_to_mem[1] ? n978 : r2[25];   // insn_decoder.v(625)
    assign n1620 = r_to_mem[1] ? n981 : r2[24];   // insn_decoder.v(625)
    assign n1621 = r_to_mem[1] ? n984 : r2[23];   // insn_decoder.v(625)
    assign n1622 = r_to_mem[1] ? n987 : r2[22];   // insn_decoder.v(625)
    assign n1623 = r_to_mem[1] ? n990 : r2[21];   // insn_decoder.v(625)
    assign n1624 = r_to_mem[1] ? n993 : r2[20];   // insn_decoder.v(625)
    assign n1625 = r_to_mem[1] ? n996 : r2[19];   // insn_decoder.v(625)
    assign n1626 = r_to_mem[1] ? n999 : r2[18];   // insn_decoder.v(625)
    assign n1627 = r_to_mem[1] ? n1002 : r2[17];   // insn_decoder.v(625)
    assign n1628 = r_to_mem[1] ? n1005 : r2[16];   // insn_decoder.v(625)
    assign n1629 = r_to_mem[1] ? n1008 : r2[15];   // insn_decoder.v(625)
    assign n1630 = r_to_mem[1] ? n1011 : r2[14];   // insn_decoder.v(625)
    assign n1631 = r_to_mem[1] ? n1014 : r2[13];   // insn_decoder.v(625)
    assign n1632 = r_to_mem[1] ? n1017 : r2[12];   // insn_decoder.v(625)
    assign n1633 = r_to_mem[1] ? n1020 : r2[11];   // insn_decoder.v(625)
    assign n1634 = r_to_mem[1] ? n1023 : r2[10];   // insn_decoder.v(625)
    assign n1635 = r_to_mem[1] ? n1026 : r2[9];   // insn_decoder.v(625)
    assign n1636 = r_to_mem[1] ? n1029 : r2[8];   // insn_decoder.v(625)
    assign n1637 = r_to_mem[1] ? n1032 : r2[7];   // insn_decoder.v(625)
    assign n1638 = r_to_mem[1] ? n1035 : r2[6];   // insn_decoder.v(625)
    assign n1639 = r_to_mem[1] ? n1038 : r2[5];   // insn_decoder.v(625)
    assign n1640 = r_to_mem[1] ? n1041 : r2[4];   // insn_decoder.v(625)
    assign n1641 = r_to_mem[1] ? n1044 : r2[3];   // insn_decoder.v(625)
    assign n1642 = r_to_mem[1] ? n1047 : r2[2];   // insn_decoder.v(625)
    assign n1643 = r_to_mem[1] ? n1050 : r2[1];   // insn_decoder.v(625)
    assign n1644 = r_to_mem[1] ? n1053 : r2[0];   // insn_decoder.v(625)
    assign n1645 = r_read[1] ? n1581 : n1225;   // insn_decoder.v(623)
    assign n1646 = r_read[1] ? n1582 : n1227;   // insn_decoder.v(623)
    assign n1647 = r_read[1] ? n1583 : n1229;   // insn_decoder.v(623)
    assign n1648 = r_read[1] ? n1584 : n1231;   // insn_decoder.v(623)
    assign n1649 = r_read[1] ? n1585 : n1233;   // insn_decoder.v(623)
    assign n1650 = r_read[1] ? n1586 : n1235;   // insn_decoder.v(623)
    assign n1651 = r_read[1] ? n1587 : n1237;   // insn_decoder.v(623)
    assign n1652 = r_read[1] ? n1588 : n1239;   // insn_decoder.v(623)
    assign n1653 = r_read[1] ? n1589 : n1241;   // insn_decoder.v(623)
    assign n1654 = r_read[1] ? n1590 : n1243;   // insn_decoder.v(623)
    assign n1655 = r_read[1] ? n1591 : n1245;   // insn_decoder.v(623)
    assign n1656 = r_read[1] ? n1592 : n1247;   // insn_decoder.v(623)
    assign n1657 = r_read[1] ? n1593 : n1249;   // insn_decoder.v(623)
    assign n1658 = r_read[1] ? n1594 : n1251;   // insn_decoder.v(623)
    assign n1659 = r_read[1] ? n1595 : n1253;   // insn_decoder.v(623)
    assign n1660 = r_read[1] ? n1596 : n1255;   // insn_decoder.v(623)
    assign n1661 = r_read[1] ? n1597 : n1257;   // insn_decoder.v(623)
    assign n1662 = r_read[1] ? n1598 : n1259;   // insn_decoder.v(623)
    assign n1663 = r_read[1] ? n1599 : n1261;   // insn_decoder.v(623)
    assign n1664 = r_read[1] ? n1600 : n1263;   // insn_decoder.v(623)
    assign n1665 = r_read[1] ? n1601 : n1265;   // insn_decoder.v(623)
    assign n1666 = r_read[1] ? n1602 : n1267;   // insn_decoder.v(623)
    assign n1667 = r_read[1] ? n1603 : n1269;   // insn_decoder.v(623)
    assign n1668 = r_read[1] ? n1604 : n1271;   // insn_decoder.v(623)
    assign n1669 = r_read[1] ? n1605 : n1273;   // insn_decoder.v(623)
    assign n1670 = r_read[1] ? n1606 : n1275;   // insn_decoder.v(623)
    assign n1671 = r_read[1] ? n1607 : n1277;   // insn_decoder.v(623)
    assign n1672 = r_read[1] ? n1608 : n1279;   // insn_decoder.v(623)
    assign n1673 = r_read[1] ? n1609 : n1281;   // insn_decoder.v(623)
    assign n1674 = r_read[1] ? n1610 : n1283;   // insn_decoder.v(623)
    assign n1675 = r_read[1] ? n1611 : n1285;   // insn_decoder.v(623)
    assign n1676 = r_read[1] ? n1612 : n1287;   // insn_decoder.v(623)
    assign n1677 = r_read[1] ? n1613 : n960;   // insn_decoder.v(623)
    assign n1678 = r_read[1] ? n1614 : n963;   // insn_decoder.v(623)
    assign n1679 = r_read[1] ? n1615 : n966;   // insn_decoder.v(623)
    assign n1680 = r_read[1] ? n1616 : n969;   // insn_decoder.v(623)
    assign n1681 = r_read[1] ? n1617 : n972;   // insn_decoder.v(623)
    assign n1682 = r_read[1] ? n1618 : n975;   // insn_decoder.v(623)
    assign n1683 = r_read[1] ? n1619 : n978;   // insn_decoder.v(623)
    assign n1684 = r_read[1] ? n1620 : n981;   // insn_decoder.v(623)
    assign n1685 = r_read[1] ? n1621 : n984;   // insn_decoder.v(623)
    assign n1686 = r_read[1] ? n1622 : n987;   // insn_decoder.v(623)
    assign n1687 = r_read[1] ? n1623 : n990;   // insn_decoder.v(623)
    assign n1688 = r_read[1] ? n1624 : n993;   // insn_decoder.v(623)
    assign n1689 = r_read[1] ? n1625 : n996;   // insn_decoder.v(623)
    assign n1690 = r_read[1] ? n1626 : n999;   // insn_decoder.v(623)
    assign n1691 = r_read[1] ? n1627 : n1002;   // insn_decoder.v(623)
    assign n1692 = r_read[1] ? n1628 : n1005;   // insn_decoder.v(623)
    assign n1693 = r_read[1] ? n1629 : n1008;   // insn_decoder.v(623)
    assign n1694 = r_read[1] ? n1630 : n1011;   // insn_decoder.v(623)
    assign n1695 = r_read[1] ? n1631 : n1014;   // insn_decoder.v(623)
    assign n1696 = r_read[1] ? n1632 : n1017;   // insn_decoder.v(623)
    assign n1697 = r_read[1] ? n1633 : n1020;   // insn_decoder.v(623)
    assign n1698 = r_read[1] ? n1634 : n1023;   // insn_decoder.v(623)
    assign n1699 = r_read[1] ? n1635 : n1026;   // insn_decoder.v(623)
    assign n1700 = r_read[1] ? n1636 : n1029;   // insn_decoder.v(623)
    assign n1701 = r_read[1] ? n1637 : n1032;   // insn_decoder.v(623)
    assign n1702 = r_read[1] ? n1638 : n1035;   // insn_decoder.v(623)
    assign n1703 = r_read[1] ? n1639 : n1038;   // insn_decoder.v(623)
    assign n1704 = r_read[1] ? n1640 : n1041;   // insn_decoder.v(623)
    assign n1705 = r_read[1] ? n1641 : n1044;   // insn_decoder.v(623)
    assign n1706 = r_read[1] ? n1642 : n1047;   // insn_decoder.v(623)
    assign n1707 = r_read[1] ? n1643 : n1050;   // insn_decoder.v(623)
    assign n1708 = r_read[1] ? n1644 : n1053;   // insn_decoder.v(623)
    assign n1709 = reg_fetch ? n1517 : n1161;   // insn_decoder.v(618)
    assign n1710 = reg_fetch ? n1518 : n1163;   // insn_decoder.v(618)
    assign n1711 = reg_fetch ? n1519 : n1165;   // insn_decoder.v(618)
    assign n1712 = reg_fetch ? n1520 : n1167;   // insn_decoder.v(618)
    assign n1713 = reg_fetch ? n1521 : n1169;   // insn_decoder.v(618)
    assign n1714 = reg_fetch ? n1522 : n1171;   // insn_decoder.v(618)
    assign n1715 = reg_fetch ? n1523 : n1173;   // insn_decoder.v(618)
    assign n1716 = reg_fetch ? n1524 : n1175;   // insn_decoder.v(618)
    assign n1717 = reg_fetch ? n1525 : n1177;   // insn_decoder.v(618)
    assign n1718 = reg_fetch ? n1526 : n1179;   // insn_decoder.v(618)
    assign n1719 = reg_fetch ? n1527 : n1181;   // insn_decoder.v(618)
    assign n1720 = reg_fetch ? n1528 : n1183;   // insn_decoder.v(618)
    assign n1721 = reg_fetch ? n1529 : n1185;   // insn_decoder.v(618)
    assign n1722 = reg_fetch ? n1530 : n1187;   // insn_decoder.v(618)
    assign n1723 = reg_fetch ? n1531 : n1189;   // insn_decoder.v(618)
    assign n1724 = reg_fetch ? n1532 : n1191;   // insn_decoder.v(618)
    assign n1725 = reg_fetch ? n1533 : n1193;   // insn_decoder.v(618)
    assign n1726 = reg_fetch ? n1534 : n1195;   // insn_decoder.v(618)
    assign n1727 = reg_fetch ? n1535 : n1197;   // insn_decoder.v(618)
    assign n1728 = reg_fetch ? n1536 : n1199;   // insn_decoder.v(618)
    assign n1729 = reg_fetch ? n1537 : n1201;   // insn_decoder.v(618)
    assign n1730 = reg_fetch ? n1538 : n1203;   // insn_decoder.v(618)
    assign n1731 = reg_fetch ? n1539 : n1205;   // insn_decoder.v(618)
    assign n1732 = reg_fetch ? n1540 : n1207;   // insn_decoder.v(618)
    assign n1733 = reg_fetch ? n1541 : n1209;   // insn_decoder.v(618)
    assign n1734 = reg_fetch ? n1542 : n1211;   // insn_decoder.v(618)
    assign n1735 = reg_fetch ? n1543 : n1213;   // insn_decoder.v(618)
    assign n1736 = reg_fetch ? n1544 : n1215;   // insn_decoder.v(618)
    assign n1737 = reg_fetch ? n1545 : n1217;   // insn_decoder.v(618)
    assign n1738 = reg_fetch ? n1546 : n1219;   // insn_decoder.v(618)
    assign n1739 = reg_fetch ? n1547 : n1221;   // insn_decoder.v(618)
    assign n1740 = reg_fetch ? n1548 : n1223;   // insn_decoder.v(618)
    assign n1741 = reg_fetch ? n1549 : n1097;   // insn_decoder.v(618)
    assign n1742 = reg_fetch ? n1550 : n1099;   // insn_decoder.v(618)
    assign n1743 = reg_fetch ? n1551 : n1101;   // insn_decoder.v(618)
    assign n1744 = reg_fetch ? n1552 : n1103;   // insn_decoder.v(618)
    assign n1745 = reg_fetch ? n1553 : n1105;   // insn_decoder.v(618)
    assign n1746 = reg_fetch ? n1554 : n1107;   // insn_decoder.v(618)
    assign n1747 = reg_fetch ? n1555 : n1109;   // insn_decoder.v(618)
    assign n1748 = reg_fetch ? n1556 : n1111;   // insn_decoder.v(618)
    assign n1749 = reg_fetch ? n1557 : n1113;   // insn_decoder.v(618)
    assign n1750 = reg_fetch ? n1558 : n1115;   // insn_decoder.v(618)
    assign n1751 = reg_fetch ? n1559 : n1117;   // insn_decoder.v(618)
    assign n1752 = reg_fetch ? n1560 : n1119;   // insn_decoder.v(618)
    assign n1753 = reg_fetch ? n1561 : n1121;   // insn_decoder.v(618)
    assign n1754 = reg_fetch ? n1562 : n1123;   // insn_decoder.v(618)
    assign n1755 = reg_fetch ? n1563 : n1125;   // insn_decoder.v(618)
    assign n1756 = reg_fetch ? n1564 : n1127;   // insn_decoder.v(618)
    assign n1757 = reg_fetch ? n1565 : n1129;   // insn_decoder.v(618)
    assign n1758 = reg_fetch ? n1566 : n1131;   // insn_decoder.v(618)
    assign n1759 = reg_fetch ? n1567 : n1133;   // insn_decoder.v(618)
    assign n1760 = reg_fetch ? n1568 : n1135;   // insn_decoder.v(618)
    assign n1761 = reg_fetch ? n1569 : n1137;   // insn_decoder.v(618)
    assign n1762 = reg_fetch ? n1570 : n1139;   // insn_decoder.v(618)
    assign n1763 = reg_fetch ? n1571 : n1141;   // insn_decoder.v(618)
    assign n1764 = reg_fetch ? n1572 : n1143;   // insn_decoder.v(618)
    assign n1765 = reg_fetch ? n1573 : n1145;   // insn_decoder.v(618)
    assign n1766 = reg_fetch ? n1574 : n1147;   // insn_decoder.v(618)
    assign n1767 = reg_fetch ? n1575 : n1149;   // insn_decoder.v(618)
    assign n1768 = reg_fetch ? n1576 : n1151;   // insn_decoder.v(618)
    assign n1769 = reg_fetch ? n1577 : n1153;   // insn_decoder.v(618)
    assign n1770 = reg_fetch ? n1578 : n1155;   // insn_decoder.v(618)
    assign n1771 = reg_fetch ? n1579 : n1157;   // insn_decoder.v(618)
    assign n1772 = reg_fetch ? n1580 : n1159;   // insn_decoder.v(618)
    assign n1773 = reg_fetch ? n1645 : n1225;   // insn_decoder.v(618)
    assign n1774 = reg_fetch ? n1646 : n1227;   // insn_decoder.v(618)
    assign n1775 = reg_fetch ? n1647 : n1229;   // insn_decoder.v(618)
    assign n1776 = reg_fetch ? n1648 : n1231;   // insn_decoder.v(618)
    assign n1777 = reg_fetch ? n1649 : n1233;   // insn_decoder.v(618)
    assign n1778 = reg_fetch ? n1650 : n1235;   // insn_decoder.v(618)
    assign n1779 = reg_fetch ? n1651 : n1237;   // insn_decoder.v(618)
    assign n1780 = reg_fetch ? n1652 : n1239;   // insn_decoder.v(618)
    assign n1781 = reg_fetch ? n1653 : n1241;   // insn_decoder.v(618)
    assign n1782 = reg_fetch ? n1654 : n1243;   // insn_decoder.v(618)
    assign n1783 = reg_fetch ? n1655 : n1245;   // insn_decoder.v(618)
    assign n1784 = reg_fetch ? n1656 : n1247;   // insn_decoder.v(618)
    assign n1785 = reg_fetch ? n1657 : n1249;   // insn_decoder.v(618)
    assign n1786 = reg_fetch ? n1658 : n1251;   // insn_decoder.v(618)
    assign n1787 = reg_fetch ? n1659 : n1253;   // insn_decoder.v(618)
    assign n1788 = reg_fetch ? n1660 : n1255;   // insn_decoder.v(618)
    assign n1789 = reg_fetch ? n1661 : n1257;   // insn_decoder.v(618)
    assign n1790 = reg_fetch ? n1662 : n1259;   // insn_decoder.v(618)
    assign n1791 = reg_fetch ? n1663 : n1261;   // insn_decoder.v(618)
    assign n1792 = reg_fetch ? n1664 : n1263;   // insn_decoder.v(618)
    assign n1793 = reg_fetch ? n1665 : n1265;   // insn_decoder.v(618)
    assign n1794 = reg_fetch ? n1666 : n1267;   // insn_decoder.v(618)
    assign n1795 = reg_fetch ? n1667 : n1269;   // insn_decoder.v(618)
    assign n1796 = reg_fetch ? n1668 : n1271;   // insn_decoder.v(618)
    assign n1797 = reg_fetch ? n1669 : n1273;   // insn_decoder.v(618)
    assign n1798 = reg_fetch ? n1670 : n1275;   // insn_decoder.v(618)
    assign n1799 = reg_fetch ? n1671 : n1277;   // insn_decoder.v(618)
    assign n1800 = reg_fetch ? n1672 : n1279;   // insn_decoder.v(618)
    assign n1801 = reg_fetch ? n1673 : n1281;   // insn_decoder.v(618)
    assign n1802 = reg_fetch ? n1674 : n1283;   // insn_decoder.v(618)
    assign n1803 = reg_fetch ? n1675 : n1285;   // insn_decoder.v(618)
    assign n1804 = reg_fetch ? n1676 : n1287;   // insn_decoder.v(618)
    assign n1805 = reg_fetch ? n1677 : n960;   // insn_decoder.v(618)
    assign n1806 = reg_fetch ? n1678 : n963;   // insn_decoder.v(618)
    assign n1807 = reg_fetch ? n1679 : n966;   // insn_decoder.v(618)
    assign n1808 = reg_fetch ? n1680 : n969;   // insn_decoder.v(618)
    assign n1809 = reg_fetch ? n1681 : n972;   // insn_decoder.v(618)
    assign n1810 = reg_fetch ? n1682 : n975;   // insn_decoder.v(618)
    assign n1811 = reg_fetch ? n1683 : n978;   // insn_decoder.v(618)
    assign n1812 = reg_fetch ? n1684 : n981;   // insn_decoder.v(618)
    assign n1813 = reg_fetch ? n1685 : n984;   // insn_decoder.v(618)
    assign n1814 = reg_fetch ? n1686 : n987;   // insn_decoder.v(618)
    assign n1815 = reg_fetch ? n1687 : n990;   // insn_decoder.v(618)
    assign n1816 = reg_fetch ? n1688 : n993;   // insn_decoder.v(618)
    assign n1817 = reg_fetch ? n1689 : n996;   // insn_decoder.v(618)
    assign n1818 = reg_fetch ? n1690 : n999;   // insn_decoder.v(618)
    assign n1819 = reg_fetch ? n1691 : n1002;   // insn_decoder.v(618)
    assign n1820 = reg_fetch ? n1692 : n1005;   // insn_decoder.v(618)
    assign n1821 = reg_fetch ? n1693 : n1008;   // insn_decoder.v(618)
    assign n1822 = reg_fetch ? n1694 : n1011;   // insn_decoder.v(618)
    assign n1823 = reg_fetch ? n1695 : n1014;   // insn_decoder.v(618)
    assign n1824 = reg_fetch ? n1696 : n1017;   // insn_decoder.v(618)
    assign n1825 = reg_fetch ? n1697 : n1020;   // insn_decoder.v(618)
    assign n1826 = reg_fetch ? n1698 : n1023;   // insn_decoder.v(618)
    assign n1827 = reg_fetch ? n1699 : n1026;   // insn_decoder.v(618)
    assign n1828 = reg_fetch ? n1700 : n1029;   // insn_decoder.v(618)
    assign n1829 = reg_fetch ? n1701 : n1032;   // insn_decoder.v(618)
    assign n1830 = reg_fetch ? n1702 : n1035;   // insn_decoder.v(618)
    assign n1831 = reg_fetch ? n1703 : n1038;   // insn_decoder.v(618)
    assign n1832 = reg_fetch ? n1704 : n1041;   // insn_decoder.v(618)
    assign n1833 = reg_fetch ? n1705 : n1044;   // insn_decoder.v(618)
    assign n1834 = reg_fetch ? n1706 : n1047;   // insn_decoder.v(618)
    assign n1835 = reg_fetch ? n1707 : n1050;   // insn_decoder.v(618)
    assign n1836 = reg_fetch ? n1708 : n1053;   // insn_decoder.v(618)
    assign n1837 = reg_fetch ? 1'b0 : n1444;   // insn_decoder.v(618)
    VERIFIC_DFFRS i1835 (.d(n1742), .clk(clk), .s(1'b0), .r(rst), .q(e_a[30]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1836 (.d(n1743), .clk(clk), .s(1'b0), .r(rst), .q(e_a[29]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1837 (.d(n1744), .clk(clk), .s(1'b0), .r(rst), .q(e_a[28]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1838 (.d(n1745), .clk(clk), .s(1'b0), .r(rst), .q(e_a[27]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1839 (.d(n1746), .clk(clk), .s(1'b0), .r(rst), .q(e_a[26]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1840 (.d(n1747), .clk(clk), .s(1'b0), .r(rst), .q(e_a[25]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1841 (.d(n1748), .clk(clk), .s(1'b0), .r(rst), .q(e_a[24]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1842 (.d(n1749), .clk(clk), .s(1'b0), .r(rst), .q(e_a[23]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1843 (.d(n1750), .clk(clk), .s(1'b0), .r(rst), .q(e_a[22]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1844 (.d(n1751), .clk(clk), .s(1'b0), .r(rst), .q(e_a[21]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1845 (.d(n1752), .clk(clk), .s(1'b0), .r(rst), .q(e_a[20]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1846 (.d(n1753), .clk(clk), .s(1'b0), .r(rst), .q(e_a[19]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1847 (.d(n1754), .clk(clk), .s(1'b0), .r(rst), .q(e_a[18]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1848 (.d(n1755), .clk(clk), .s(1'b0), .r(rst), .q(e_a[17]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1849 (.d(n1756), .clk(clk), .s(1'b0), .r(rst), .q(e_a[16]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1850 (.d(n1757), .clk(clk), .s(1'b0), .r(rst), .q(e_a[15]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1851 (.d(n1758), .clk(clk), .s(1'b0), .r(rst), .q(e_a[14]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1852 (.d(n1759), .clk(clk), .s(1'b0), .r(rst), .q(e_a[13]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1853 (.d(n1760), .clk(clk), .s(1'b0), .r(rst), .q(e_a[12]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1854 (.d(n1761), .clk(clk), .s(1'b0), .r(rst), .q(e_a[11]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1855 (.d(n1762), .clk(clk), .s(1'b0), .r(rst), .q(e_a[10]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1856 (.d(n1763), .clk(clk), .s(1'b0), .r(rst), .q(e_a[9]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1857 (.d(n1764), .clk(clk), .s(1'b0), .r(rst), .q(e_a[8]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1858 (.d(n1765), .clk(clk), .s(1'b0), .r(rst), .q(e_a[7]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1859 (.d(n1766), .clk(clk), .s(1'b0), .r(rst), .q(e_a[6]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1860 (.d(n1767), .clk(clk), .s(1'b0), .r(rst), .q(e_a[5]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1861 (.d(n1768), .clk(clk), .s(1'b0), .r(rst), .q(e_a[4]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1862 (.d(n1769), .clk(clk), .s(1'b0), .r(rst), .q(e_a[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1863 (.d(n1770), .clk(clk), .s(1'b0), .r(rst), .q(e_a[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1864 (.d(n1771), .clk(clk), .s(1'b0), .r(rst), .q(e_a[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1865 (.d(n1772), .clk(clk), .s(1'b0), .r(rst), .q(e_a[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1866 (.d(n1805), .clk(clk), .s(1'b0), .r(rst), .q(e_b[31]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1867 (.d(n1806), .clk(clk), .s(1'b0), .r(rst), .q(e_b[30]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1868 (.d(n1807), .clk(clk), .s(1'b0), .r(rst), .q(e_b[29]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1869 (.d(n1808), .clk(clk), .s(1'b0), .r(rst), .q(e_b[28]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1870 (.d(n1809), .clk(clk), .s(1'b0), .r(rst), .q(e_b[27]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1871 (.d(n1810), .clk(clk), .s(1'b0), .r(rst), .q(e_b[26]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1872 (.d(n1811), .clk(clk), .s(1'b0), .r(rst), .q(e_b[25]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1873 (.d(n1812), .clk(clk), .s(1'b0), .r(rst), .q(e_b[24]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1874 (.d(n1813), .clk(clk), .s(1'b0), .r(rst), .q(e_b[23]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1875 (.d(n1814), .clk(clk), .s(1'b0), .r(rst), .q(e_b[22]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1876 (.d(n1815), .clk(clk), .s(1'b0), .r(rst), .q(e_b[21]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1877 (.d(n1816), .clk(clk), .s(1'b0), .r(rst), .q(e_b[20]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1878 (.d(n1817), .clk(clk), .s(1'b0), .r(rst), .q(e_b[19]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1879 (.d(n1818), .clk(clk), .s(1'b0), .r(rst), .q(e_b[18]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1880 (.d(n1819), .clk(clk), .s(1'b0), .r(rst), .q(e_b[17]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1881 (.d(n1820), .clk(clk), .s(1'b0), .r(rst), .q(e_b[16]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1882 (.d(n1821), .clk(clk), .s(1'b0), .r(rst), .q(e_b[15]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1883 (.d(n1822), .clk(clk), .s(1'b0), .r(rst), .q(e_b[14]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1884 (.d(n1823), .clk(clk), .s(1'b0), .r(rst), .q(e_b[13]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1885 (.d(n1824), .clk(clk), .s(1'b0), .r(rst), .q(e_b[12]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1886 (.d(n1825), .clk(clk), .s(1'b0), .r(rst), .q(e_b[11]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1887 (.d(n1826), .clk(clk), .s(1'b0), .r(rst), .q(e_b[10]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1888 (.d(n1827), .clk(clk), .s(1'b0), .r(rst), .q(e_b[9]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1889 (.d(n1828), .clk(clk), .s(1'b0), .r(rst), .q(e_b[8]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1890 (.d(n1829), .clk(clk), .s(1'b0), .r(rst), .q(e_b[7]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1891 (.d(n1830), .clk(clk), .s(1'b0), .r(rst), .q(e_b[6]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1892 (.d(n1831), .clk(clk), .s(1'b0), .r(rst), .q(e_b[5]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1893 (.d(n1832), .clk(clk), .s(1'b0), .r(rst), .q(e_b[4]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1894 (.d(n1833), .clk(clk), .s(1'b0), .r(rst), .q(e_b[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1895 (.d(n1834), .clk(clk), .s(1'b0), .r(rst), .q(e_b[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1896 (.d(n1835), .clk(clk), .s(1'b0), .r(rst), .q(e_b[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1897 (.d(n1836), .clk(clk), .s(1'b0), .r(rst), .q(e_b[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1898 (.d(n772), .clk(clk), .s(1'b0), .r(rst), .q(e_alu_op[7]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1899 (.d(n774), .clk(clk), .s(1'b0), .r(rst), .q(e_alu_op[6]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1900 (.d(n776), .clk(clk), .s(1'b0), .r(rst), .q(e_alu_op[5]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1901 (.d(n780), .clk(clk), .s(1'b0), .r(rst), .q(e_alu_op[4]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1902 (.d(n784), .clk(clk), .s(1'b0), .r(rst), .q(e_alu_op[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1903 (.d(n788), .clk(clk), .s(1'b0), .r(rst), .q(e_alu_op[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1904 (.d(n792), .clk(clk), .s(1'b0), .r(rst), .q(e_alu_op[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1905 (.d(n796), .clk(clk), .s(1'b0), .r(rst), .q(e_alu_op[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1906 (.d(n799), .clk(clk), .s(1'b0), .r(rst), .q(e_cond[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1907 (.d(n802), .clk(clk), .s(1'b0), .r(rst), .q(e_cond[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1908 (.d(n805), .clk(clk), .s(1'b0), .r(rst), .q(e_cond[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1909 (.d(n808), .clk(clk), .s(1'b0), .r(rst), .q(e_cond[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1910 (.d(n812), .clk(clk), .s(1'b0), .r(rst), .q(e_write_flags[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1911 (.d(n816), .clk(clk), .s(1'b0), .r(rst), .q(e_write_flags[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1912 (.d(n820), .clk(clk), .s(1'b0), .r(rst), .q(e_write_flags[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1913 (.d(n824), .clk(clk), .s(1'b0), .r(rst), .q(e_write_flags[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1914 (.d(e_swp), .clk(clk), .s(1'b0), .r(rst), .q(e_swp));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1915 (.d(n827), .clk(clk), .s(1'b0), .r(rst), .q(e_is_cond));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1916 (.d(n1709), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[31]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1917 (.d(n1710), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[30]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1918 (.d(n1711), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[29]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1919 (.d(n1712), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[28]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1920 (.d(n1713), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[27]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1921 (.d(n1714), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[26]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1922 (.d(n1715), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[25]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1923 (.d(n1716), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[24]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1924 (.d(n1717), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[23]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1925 (.d(n1718), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[22]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1926 (.d(n1719), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[21]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1927 (.d(n1720), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[20]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1928 (.d(n1721), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[19]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1929 (.d(n1722), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[18]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1930 (.d(n1723), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[17]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1931 (.d(n1724), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[16]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1932 (.d(n1725), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[15]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1933 (.d(n1726), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[14]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1934 (.d(n1727), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[13]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1935 (.d(n1728), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[12]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1936 (.d(n1729), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[11]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1937 (.d(n1730), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[10]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1938 (.d(n1731), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[9]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1939 (.d(n1732), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[8]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1940 (.d(n1733), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[7]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1941 (.d(n1734), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[6]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1942 (.d(n1735), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[5]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1943 (.d(n1736), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[4]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1944 (.d(n1737), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1945 (.d(n1738), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1946 (.d(n1739), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1947 (.d(n1740), .clk(clk), .s(1'b0), .r(rst), .q(m_a1[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1948 (.d(n1773), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[31]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1949 (.d(n1774), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[30]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1950 (.d(n1775), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[29]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1951 (.d(n1776), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[28]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1952 (.d(n1777), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[27]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1953 (.d(n1778), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[26]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1954 (.d(n1779), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[25]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1955 (.d(n1780), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[24]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1956 (.d(n1781), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[23]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1957 (.d(n1782), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[22]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1958 (.d(n1783), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[21]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1959 (.d(n1784), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[20]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1960 (.d(n1785), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[19]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1961 (.d(n1786), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[18]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1962 (.d(n1787), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[17]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1963 (.d(n1788), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[16]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1964 (.d(n1789), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[15]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1965 (.d(n1790), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[14]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1966 (.d(n1791), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[13]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1967 (.d(n1792), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[12]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1968 (.d(n1793), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[11]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1969 (.d(n1794), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[10]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1970 (.d(n1795), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[9]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1971 (.d(n1796), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[8]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1972 (.d(n1797), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[7]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1973 (.d(n1798), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[6]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1974 (.d(n1799), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[5]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1975 (.d(n1800), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[4]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1976 (.d(n1801), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1977 (.d(n1802), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1978 (.d(n1803), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1979 (.d(n1804), .clk(clk), .s(1'b0), .r(rst), .q(m_a2[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1980 (.d(n830), .clk(clk), .s(1'b0), .r(rst), .q(m_r1_op[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1981 (.d(n832), .clk(clk), .s(1'b0), .r(rst), .q(m_r1_op[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1982 (.d(n835), .clk(clk), .s(1'b0), .r(rst), .q(m_r1_op[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1983 (.d(n839), .clk(clk), .s(1'b0), .r(rst), .q(m_r1_op[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1984 (.d(n842), .clk(clk), .s(1'b0), .r(rst), .q(m_r2_op[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1985 (.d(n845), .clk(clk), .s(1'b0), .r(rst), .q(m_r2_op[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1986 (.d(n848), .clk(clk), .s(1'b0), .r(rst), .q(m_r2_op[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1987 (.d(n851), .clk(clk), .s(1'b0), .r(rst), .q(m_r2_op[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1988 (.d(n882), .clk(clk), .s(1'b0), .r(rst), .q(r_a1[4]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1989 (.d(n886), .clk(clk), .s(1'b0), .r(rst), .q(r_a1[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1990 (.d(n890), .clk(clk), .s(1'b0), .r(rst), .q(r_a1[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1991 (.d(n894), .clk(clk), .s(1'b0), .r(rst), .q(r_a1[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1992 (.d(n898), .clk(clk), .s(1'b0), .r(rst), .q(r_a1[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1993 (.d(n945), .clk(clk), .s(1'b0), .r(rst), .q(r_a2[4]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1994 (.d(n948), .clk(clk), .s(1'b0), .r(rst), .q(r_a2[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1995 (.d(n951), .clk(clk), .s(1'b0), .r(rst), .q(r_a2[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1996 (.d(n954), .clk(clk), .s(1'b0), .r(rst), .q(r_a2[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1997 (.d(n957), .clk(clk), .s(1'b0), .r(rst), .q(r_a2[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1998 (.d(n853), .clk(clk), .s(1'b0), .r(rst), .q(r_op[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i1999 (.d(n857), .clk(clk), .s(1'b0), .r(rst), .q(r_op[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2000 (.d(n861), .clk(clk), .s(1'b0), .r(rst), .q(r_op[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2001 (.d(n865), .clk(clk), .s(1'b0), .r(rst), .q(r_op[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2002 (.d(n1442), .clk(clk), .s(1'b0), .r(rst), .q(d_pass));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2004 (.d(n902), .clk(clk), .s(1'b0), .r(rst), .q(r_r1_addr[4]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2005 (.d(n906), .clk(clk), .s(1'b0), .r(rst), .q(r_r1_addr[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2006 (.d(n910), .clk(clk), .s(1'b0), .r(rst), .q(r_r1_addr[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2007 (.d(n913), .clk(clk), .s(1'b0), .r(rst), .q(r_r1_addr[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2008 (.d(n917), .clk(clk), .s(1'b0), .r(rst), .q(r_r1_addr[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2009 (.d(n920), .clk(clk), .s(1'b0), .r(rst), .q(r_r2_addr[4]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2010 (.d(n923), .clk(clk), .s(1'b0), .r(rst), .q(r_r2_addr[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2011 (.d(n926), .clk(clk), .s(1'b0), .r(rst), .q(r_r2_addr[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2012 (.d(n929), .clk(clk), .s(1'b0), .r(rst), .q(r_r2_addr[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2013 (.d(n932), .clk(clk), .s(1'b0), .r(rst), .q(r_r2_addr[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2014 (.d(n1401), .clk(clk), .s(1'b0), .r(rst), .q(r_read[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2015 (.d(n1402), .clk(clk), .s(1'b0), .r(rst), .q(r_read[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2016 (.d(n1445), .clk(clk), .s(1'b0), .r(rst), .q(state1[7]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2017 (.d(n1446), .clk(clk), .s(1'b0), .r(rst), .q(state1[6]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2018 (.d(n1447), .clk(clk), .s(1'b0), .r(rst), .q(state1[5]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2019 (.d(n1448), .clk(clk), .s(1'b0), .r(rst), .q(state1[4]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2020 (.d(n1449), .clk(clk), .s(1'b0), .r(rst), .q(state1[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2021 (.d(n1450), .clk(clk), .s(1'b0), .r(rst), .q(state1[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2022 (.d(n1451), .clk(clk), .s(1'b0), .r(rst), .q(state1[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2023 (.d(n1452), .clk(clk), .s(1'b0), .r(rst), .q(state1[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2024 (.d(n1443), .clk(clk), .s(rst), .r(1'b0), .q(fetch));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2025 (.d(n1837), .clk(clk), .s(1'b0), .r(rst), .q(reg_fetch));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2026 (.d(n1411), .clk(clk), .s(1'b0), .r(rst), .q(old_pass_imm));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2027 (.d(n1412), .clk(clk), .s(1'b0), .r(rst), .q(old_fetch_imm));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2028 (.d(n1413), .clk(clk), .s(1'b0), .r(rst), .q(old_pcincr_imm));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2029 (.d(n1403), .clk(clk), .s(1'b0), .r(rst), .q(old_state1_imm[7]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2030 (.d(n1404), .clk(clk), .s(1'b0), .r(rst), .q(old_state1_imm[6]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2031 (.d(n1405), .clk(clk), .s(1'b0), .r(rst), .q(old_state1_imm[5]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2032 (.d(n1406), .clk(clk), .s(1'b0), .r(rst), .q(old_state1_imm[4]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2033 (.d(n1407), .clk(clk), .s(1'b0), .r(rst), .q(old_state1_imm[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2034 (.d(n1408), .clk(clk), .s(1'b0), .r(rst), .q(old_state1_imm[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2035 (.d(n1409), .clk(clk), .s(1'b0), .r(rst), .q(old_state1_imm[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2036 (.d(n1410), .clk(clk), .s(1'b0), .r(rst), .q(old_state1_imm[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2037 (.d(n1431), .clk(clk), .s(1'b0), .r(rst), .q(old_pass_hz));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2038 (.d(n1432), .clk(clk), .s(1'b0), .r(rst), .q(old_fetch_hz));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2039 (.d(n1430), .clk(clk), .s(1'b0), .r(rst), .q(old_pcincr_hz));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2040 (.d(n1433), .clk(clk), .s(1'b0), .r(rst), .q(old_state1_hz[7]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2041 (.d(n1434), .clk(clk), .s(1'b0), .r(rst), .q(old_state1_hz[6]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2042 (.d(n1435), .clk(clk), .s(1'b0), .r(rst), .q(old_state1_hz[5]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2043 (.d(n1436), .clk(clk), .s(1'b0), .r(rst), .q(old_state1_hz[4]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2044 (.d(n1437), .clk(clk), .s(1'b0), .r(rst), .q(old_state1_hz[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2045 (.d(n1438), .clk(clk), .s(1'b0), .r(rst), .q(old_state1_hz[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2046 (.d(n1439), .clk(clk), .s(1'b0), .r(rst), .q(old_state1_hz[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2047 (.d(n1440), .clk(clk), .s(1'b0), .r(rst), .q(old_state1_hz[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2048 (.d(n1302), .clk(clk), .s(1'b0), .r(rst), .q(set_delay));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2056 (.d(n1086), .clk(clk), .s(1'b0), .r(rst), .q(delay_counter[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2057 (.d(n1089), .clk(clk), .s(1'b0), .r(rst), .q(delay_counter[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2058 (.d(n1092), .clk(clk), .s(1'b0), .r(rst), .q(delay_counter[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2059 (.d(n1095), .clk(clk), .s(1'b0), .r(rst), .q(delay_counter[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2060 (.d(n1426), .clk(clk), .s(1'b0), .r(rst), .q(imm_action[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2061 (.d(n1427), .clk(clk), .s(1'b0), .r(rst), .q(imm_action[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2062 (.d(n1428), .clk(clk), .s(1'b0), .r(rst), .q(imm_action[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2063 (.d(n874), .clk(clk), .s(1'b0), .r(rst), .q(r_to_mem[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2064 (.d(n878), .clk(clk), .s(1'b0), .r(rst), .q(r_to_mem[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2065 (.d(n2073), .clk(clk), .s(1'b0), .r(1'b0), .q(cond[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2066 (.d(n2074), .clk(clk), .s(1'b0), .r(1'b0), .q(cond[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2067 (.d(n2075), .clk(clk), .s(1'b0), .r(1'b0), .q(cond[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2068 (.d(n2076), .clk(clk), .s(1'b0), .r(1'b0), .q(cond[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2073 (.d(n2082), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_a_addr[4]));   // insn_decoder.v(158)
    assign n2073 = rst ? cond[3] : n12;   // insn_decoder.v(158)
    assign n2074 = rst ? cond[2] : n13;   // insn_decoder.v(158)
    assign n2075 = rst ? cond[1] : n14;   // insn_decoder.v(158)
    assign n2076 = rst ? cond[0] : n15;   // insn_decoder.v(158)
    VERIFIC_DFFRS i2074 (.d(n2083), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_a_addr[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2075 (.d(n2084), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_a_addr[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2076 (.d(n2085), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_a_addr[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2077 (.d(n2086), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_a_addr[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2083 (.d(n2092), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_b_addr[4]));   // insn_decoder.v(158)
    assign n2082 = rst ? reg_a_addr[4] : n16;   // insn_decoder.v(158)
    assign n2083 = rst ? reg_a_addr[3] : n17;   // insn_decoder.v(158)
    assign n2084 = rst ? reg_a_addr[2] : n18;   // insn_decoder.v(158)
    assign n2085 = rst ? reg_a_addr[1] : n19;   // insn_decoder.v(158)
    assign n2086 = rst ? reg_a_addr[0] : n20;   // insn_decoder.v(158)
    VERIFIC_DFFRS i2084 (.d(n2093), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_b_addr[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2085 (.d(n2094), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_b_addr[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2086 (.d(n2095), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_b_addr[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2087 (.d(n2096), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_b_addr[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2093 (.d(n2102), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_c_addr[4]));   // insn_decoder.v(158)
    assign n2092 = rst ? reg_b_addr[4] : n21;   // insn_decoder.v(158)
    assign n2093 = rst ? reg_b_addr[3] : n22;   // insn_decoder.v(158)
    assign n2094 = rst ? reg_b_addr[2] : n23;   // insn_decoder.v(158)
    assign n2095 = rst ? reg_b_addr[1] : n24;   // insn_decoder.v(158)
    assign n2096 = rst ? reg_b_addr[0] : n25;   // insn_decoder.v(158)
    VERIFIC_DFFRS i2094 (.d(n2103), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_c_addr[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2095 (.d(n2104), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_c_addr[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2096 (.d(n2105), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_c_addr[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2097 (.d(n2106), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_c_addr[0]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2103 (.d(n2112), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_d_addr[4]));   // insn_decoder.v(158)
    assign n2102 = rst ? reg_c_addr[4] : n26;   // insn_decoder.v(158)
    assign n2103 = rst ? reg_c_addr[3] : n27;   // insn_decoder.v(158)
    assign n2104 = rst ? reg_c_addr[2] : n28;   // insn_decoder.v(158)
    assign n2105 = rst ? reg_c_addr[1] : n29;   // insn_decoder.v(158)
    assign n2106 = rst ? reg_c_addr[0] : n30;   // insn_decoder.v(158)
    VERIFIC_DFFRS i2104 (.d(n2113), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_d_addr[3]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2105 (.d(n2114), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_d_addr[2]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2106 (.d(n2115), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_d_addr[1]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2107 (.d(n2116), .clk(clk), .s(1'b0), .r(1'b0), .q(reg_d_addr[0]));   // insn_decoder.v(158)
    assign n2112 = rst ? reg_d_addr[4] : n31;   // insn_decoder.v(158)
    assign n2113 = rst ? reg_d_addr[3] : n32;   // insn_decoder.v(158)
    assign n2114 = rst ? reg_d_addr[2] : n33;   // insn_decoder.v(158)
    assign n2115 = rst ? reg_d_addr[1] : n34;   // insn_decoder.v(158)
    assign n2116 = rst ? reg_d_addr[0] : n35;   // insn_decoder.v(158)
    VERIFIC_DFFRS i1834 (.d(n1741), .clk(clk), .s(1'b0), .r(rst), .q(e_a[31]));   // insn_decoder.v(158)
    VERIFIC_DFFRS i2003 (.d(n1441), .clk(clk), .s(rst), .r(1'b0), .q(d_pcincr));   // insn_decoder.v(158)
    
endmodule

//
// Verific Verilog Description of OPERATOR LessThan_4u_4u
//

module LessThan_4u_4u (cin, a, b, o);
    input cin;
    input [3:0]a;
    input [3:0]b;
    output o;
    assign o = cin ? a<=b : a<b ;
    
endmodule

//
// Verific Verilog Description of OPERATOR add_4u_4u
//

module add_4u_4u (cin, a, b, o, cout);
    input cin;
    input [3:0]a;
    input [3:0]b;
    output [3:0]o;
    output cout;
    assign {cout, o} = a + b + cin;
    
endmodule

//
// Verific Verilog Description of OPERATOR Select_3
//

module Select_3 (sel, data, o);
    input [2:0]sel;
    input [2:0]data;
    output o;
    assign o = |(sel & data);
    
endmodule

//
// Verific Verilog Description of OPERATOR Select_4
//

module Select_4 (sel, data, o);
    input [3:0]sel;
    input [3:0]data;
    output o;
    assign o = |(sel & data);
    
endmodule

//
// Verific Verilog Description of OPERATOR Select_5
//

module Select_5 (sel, data, o);
    input [4:0]sel;
    input [4:0]data;
    output o;
    assign o = |(sel & data);
    
endmodule

//
// Verific Verilog Description of module pipeline_interface
//

module pipeline_interface (qe_a, qe_b, qe_alu_op, qe_is_cond, qe_cond, 
            qe_write_flags, qe_swp, qm_a1, qm_a2, qm_r1_op, qm_r2_op, 
            qr_a1, qr_a2, qr_op, qd_pcincr, e_a, e_b, e_alu_op, 
            e_is_cond, e_cond, e_write_flags, e_swp, m_a1, m_a2, 
            m_r1_op, m_r2_op, r_a1, r_a2, r_op, d_pass, d_pcincr, 
            clk, rst);   // pipeline_interface.v(3)
    output [31:0]qe_a;   // pipeline_interface.v(24)
    output [31:0]qe_b;   // pipeline_interface.v(24)
    output [7:0]qe_alu_op;   // pipeline_interface.v(25)
    output qe_is_cond;   // pipeline_interface.v(29)
    output [3:0]qe_cond;   // pipeline_interface.v(26)
    output [3:0]qe_write_flags;   // pipeline_interface.v(27)
    output qe_swp;   // pipeline_interface.v(28)
    output [31:0]qm_a1;   // pipeline_interface.v(31)
    output [31:0]qm_a2;   // pipeline_interface.v(31)
    output [3:0]qm_r1_op;   // pipeline_interface.v(32)
    output [3:0]qm_r2_op;   // pipeline_interface.v(32)
    output [4:0]qr_a1;   // pipeline_interface.v(34)
    output [4:0]qr_a2;   // pipeline_interface.v(34)
    output [3:0]qr_op;   // pipeline_interface.v(35)
    output qd_pcincr;   // pipeline_interface.v(37)
    input [31:0]e_a;   // pipeline_interface.v(6)
    input [31:0]e_b;   // pipeline_interface.v(6)
    input [7:0]e_alu_op;   // pipeline_interface.v(7)
    input e_is_cond;   // pipeline_interface.v(11)
    input [3:0]e_cond;   // pipeline_interface.v(8)
    input [3:0]e_write_flags;   // pipeline_interface.v(9)
    input e_swp;   // pipeline_interface.v(10)
    input [31:0]m_a1;   // pipeline_interface.v(13)
    input [31:0]m_a2;   // pipeline_interface.v(13)
    input [3:0]m_r1_op;   // pipeline_interface.v(14)
    input [3:0]m_r2_op;   // pipeline_interface.v(14)
    input [4:0]r_a1;   // pipeline_interface.v(16)
    input [4:0]r_a2;   // pipeline_interface.v(16)
    input [3:0]r_op;   // pipeline_interface.v(17)
    input d_pass;   // pipeline_interface.v(19)
    input d_pcincr;   // pipeline_interface.v(20)
    input clk;   // pipeline_interface.v(22)
    input rst;   // pipeline_interface.v(22)
    
    
    wire n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
        n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, 
        n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, 
        n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
        n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, 
        n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
        n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
        n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, 
        n97, n98, n99, n100, n101, n102, n103, n104, n105, 
        n106, n107, n108, n109, n110, n111, n112, n113, n114, 
        n115, n116, n117, n118, n119, n120, n121, n122, n123, 
        n124, n125, n126, n127, n128, n129, n130, n131, n132, 
        n133, n134, n135, n136, n137, n138, n139, n140, n141, 
        n142, n143, n144, n145, n146, n147, n148, n149, n150, 
        n151, n152, n153, n154, n155, n156, n157, n158, n159, 
        n160, n161, n162, n163, n164, n165, n166, n167, n168, 
        n169, n170, n171, n172, n173, n174, n175;
    
    not (n6, d_pass) ;   // pipeline_interface.v(64)
    assign n8 = n6 ? 1'b0 : e_a[31];   // pipeline_interface.v(78)
    assign n9 = n6 ? 1'b0 : e_a[30];   // pipeline_interface.v(78)
    assign n10 = n6 ? 1'b0 : e_a[29];   // pipeline_interface.v(78)
    assign n11 = n6 ? 1'b0 : e_a[28];   // pipeline_interface.v(78)
    assign n12 = n6 ? 1'b0 : e_a[27];   // pipeline_interface.v(78)
    assign n13 = n6 ? 1'b0 : e_a[26];   // pipeline_interface.v(78)
    assign n14 = n6 ? 1'b0 : e_a[25];   // pipeline_interface.v(78)
    assign n15 = n6 ? 1'b0 : e_a[24];   // pipeline_interface.v(78)
    assign n16 = n6 ? 1'b0 : e_a[23];   // pipeline_interface.v(78)
    assign n17 = n6 ? 1'b0 : e_a[22];   // pipeline_interface.v(78)
    assign n18 = n6 ? 1'b0 : e_a[21];   // pipeline_interface.v(78)
    assign n19 = n6 ? 1'b0 : e_a[20];   // pipeline_interface.v(78)
    assign n20 = n6 ? 1'b0 : e_a[19];   // pipeline_interface.v(78)
    assign n21 = n6 ? 1'b0 : e_a[18];   // pipeline_interface.v(78)
    assign n22 = n6 ? 1'b0 : e_a[17];   // pipeline_interface.v(78)
    assign n23 = n6 ? 1'b0 : e_a[16];   // pipeline_interface.v(78)
    assign n24 = n6 ? 1'b0 : e_a[15];   // pipeline_interface.v(78)
    assign n25 = n6 ? 1'b0 : e_a[14];   // pipeline_interface.v(78)
    assign n26 = n6 ? 1'b0 : e_a[13];   // pipeline_interface.v(78)
    assign n27 = n6 ? 1'b0 : e_a[12];   // pipeline_interface.v(78)
    assign n28 = n6 ? 1'b0 : e_a[11];   // pipeline_interface.v(78)
    assign n29 = n6 ? 1'b0 : e_a[10];   // pipeline_interface.v(78)
    assign n30 = n6 ? 1'b0 : e_a[9];   // pipeline_interface.v(78)
    assign n31 = n6 ? 1'b0 : e_a[8];   // pipeline_interface.v(78)
    assign n32 = n6 ? 1'b0 : e_a[7];   // pipeline_interface.v(78)
    assign n33 = n6 ? 1'b0 : e_a[6];   // pipeline_interface.v(78)
    assign n34 = n6 ? 1'b0 : e_a[5];   // pipeline_interface.v(78)
    assign n35 = n6 ? 1'b0 : e_a[4];   // pipeline_interface.v(78)
    assign n36 = n6 ? 1'b0 : e_a[3];   // pipeline_interface.v(78)
    assign n37 = n6 ? 1'b0 : e_a[2];   // pipeline_interface.v(78)
    assign n38 = n6 ? 1'b0 : e_a[1];   // pipeline_interface.v(78)
    assign n39 = n6 ? 1'b0 : e_a[0];   // pipeline_interface.v(78)
    assign n40 = n6 ? 1'b0 : e_b[31];   // pipeline_interface.v(78)
    assign n41 = n6 ? 1'b0 : e_b[30];   // pipeline_interface.v(78)
    assign n42 = n6 ? 1'b0 : e_b[29];   // pipeline_interface.v(78)
    assign n43 = n6 ? 1'b0 : e_b[28];   // pipeline_interface.v(78)
    assign n44 = n6 ? 1'b0 : e_b[27];   // pipeline_interface.v(78)
    assign n45 = n6 ? 1'b0 : e_b[26];   // pipeline_interface.v(78)
    assign n46 = n6 ? 1'b0 : e_b[25];   // pipeline_interface.v(78)
    assign n47 = n6 ? 1'b0 : e_b[24];   // pipeline_interface.v(78)
    assign n48 = n6 ? 1'b0 : e_b[23];   // pipeline_interface.v(78)
    assign n49 = n6 ? 1'b0 : e_b[22];   // pipeline_interface.v(78)
    assign n50 = n6 ? 1'b0 : e_b[21];   // pipeline_interface.v(78)
    assign n51 = n6 ? 1'b0 : e_b[20];   // pipeline_interface.v(78)
    assign n52 = n6 ? 1'b0 : e_b[19];   // pipeline_interface.v(78)
    assign n53 = n6 ? 1'b0 : e_b[18];   // pipeline_interface.v(78)
    assign n54 = n6 ? 1'b0 : e_b[17];   // pipeline_interface.v(78)
    assign n55 = n6 ? 1'b0 : e_b[16];   // pipeline_interface.v(78)
    assign n56 = n6 ? 1'b0 : e_b[15];   // pipeline_interface.v(78)
    assign n57 = n6 ? 1'b0 : e_b[14];   // pipeline_interface.v(78)
    assign n58 = n6 ? 1'b0 : e_b[13];   // pipeline_interface.v(78)
    assign n59 = n6 ? 1'b0 : e_b[12];   // pipeline_interface.v(78)
    assign n60 = n6 ? 1'b0 : e_b[11];   // pipeline_interface.v(78)
    assign n61 = n6 ? 1'b0 : e_b[10];   // pipeline_interface.v(78)
    assign n62 = n6 ? 1'b0 : e_b[9];   // pipeline_interface.v(78)
    assign n63 = n6 ? 1'b0 : e_b[8];   // pipeline_interface.v(78)
    assign n64 = n6 ? 1'b0 : e_b[7];   // pipeline_interface.v(78)
    assign n65 = n6 ? 1'b0 : e_b[6];   // pipeline_interface.v(78)
    assign n66 = n6 ? 1'b0 : e_b[5];   // pipeline_interface.v(78)
    assign n67 = n6 ? 1'b0 : e_b[4];   // pipeline_interface.v(78)
    assign n68 = n6 ? 1'b0 : e_b[3];   // pipeline_interface.v(78)
    assign n69 = n6 ? 1'b0 : e_b[2];   // pipeline_interface.v(78)
    assign n70 = n6 ? 1'b0 : e_b[1];   // pipeline_interface.v(78)
    assign n71 = n6 ? 1'b0 : e_b[0];   // pipeline_interface.v(78)
    assign n72 = n6 ? 1'b0 : e_alu_op[7];   // pipeline_interface.v(78)
    assign n73 = n6 ? 1'b0 : e_alu_op[6];   // pipeline_interface.v(78)
    assign n74 = n6 ? 1'b0 : e_alu_op[5];   // pipeline_interface.v(78)
    assign n75 = n6 ? 1'b0 : e_alu_op[4];   // pipeline_interface.v(78)
    assign n76 = n6 ? 1'b0 : e_alu_op[3];   // pipeline_interface.v(78)
    assign n77 = n6 ? 1'b0 : e_alu_op[2];   // pipeline_interface.v(78)
    assign n78 = n6 ? 1'b0 : e_alu_op[1];   // pipeline_interface.v(78)
    assign n79 = n6 ? 1'b0 : e_alu_op[0];   // pipeline_interface.v(78)
    assign n80 = n6 ? 1'b0 : e_cond[3];   // pipeline_interface.v(78)
    assign n81 = n6 ? 1'b0 : e_cond[2];   // pipeline_interface.v(78)
    assign n82 = n6 ? 1'b0 : e_cond[1];   // pipeline_interface.v(78)
    assign n83 = n6 ? 1'b0 : e_cond[0];   // pipeline_interface.v(78)
    assign n84 = n6 ? 1'b0 : e_write_flags[3];   // pipeline_interface.v(78)
    assign n85 = n6 ? 1'b0 : e_write_flags[2];   // pipeline_interface.v(78)
    assign n86 = n6 ? 1'b0 : e_write_flags[1];   // pipeline_interface.v(78)
    assign n87 = n6 ? 1'b0 : e_write_flags[0];   // pipeline_interface.v(78)
    assign n88 = n6 ? 1'b0 : e_swp;   // pipeline_interface.v(78)
    assign n89 = n6 ? 1'b0 : e_is_cond;   // pipeline_interface.v(78)
    assign n90 = n6 ? 1'b0 : m_a1[31];   // pipeline_interface.v(78)
    assign n91 = n6 ? 1'b0 : m_a1[30];   // pipeline_interface.v(78)
    assign n92 = n6 ? 1'b0 : m_a1[29];   // pipeline_interface.v(78)
    assign n93 = n6 ? 1'b0 : m_a1[28];   // pipeline_interface.v(78)
    assign n94 = n6 ? 1'b0 : m_a1[27];   // pipeline_interface.v(78)
    assign n95 = n6 ? 1'b0 : m_a1[26];   // pipeline_interface.v(78)
    assign n96 = n6 ? 1'b0 : m_a1[25];   // pipeline_interface.v(78)
    assign n97 = n6 ? 1'b0 : m_a1[24];   // pipeline_interface.v(78)
    assign n98 = n6 ? 1'b0 : m_a1[23];   // pipeline_interface.v(78)
    assign n99 = n6 ? 1'b0 : m_a1[22];   // pipeline_interface.v(78)
    assign n100 = n6 ? 1'b0 : m_a1[21];   // pipeline_interface.v(78)
    assign n101 = n6 ? 1'b0 : m_a1[20];   // pipeline_interface.v(78)
    assign n102 = n6 ? 1'b0 : m_a1[19];   // pipeline_interface.v(78)
    assign n103 = n6 ? 1'b0 : m_a1[18];   // pipeline_interface.v(78)
    assign n104 = n6 ? 1'b0 : m_a1[17];   // pipeline_interface.v(78)
    assign n105 = n6 ? 1'b0 : m_a1[16];   // pipeline_interface.v(78)
    assign n106 = n6 ? 1'b0 : m_a1[15];   // pipeline_interface.v(78)
    assign n107 = n6 ? 1'b0 : m_a1[14];   // pipeline_interface.v(78)
    assign n108 = n6 ? 1'b0 : m_a1[13];   // pipeline_interface.v(78)
    assign n109 = n6 ? 1'b0 : m_a1[12];   // pipeline_interface.v(78)
    assign n110 = n6 ? 1'b0 : m_a1[11];   // pipeline_interface.v(78)
    assign n111 = n6 ? 1'b0 : m_a1[10];   // pipeline_interface.v(78)
    assign n112 = n6 ? 1'b0 : m_a1[9];   // pipeline_interface.v(78)
    assign n113 = n6 ? 1'b0 : m_a1[8];   // pipeline_interface.v(78)
    assign n114 = n6 ? 1'b0 : m_a1[7];   // pipeline_interface.v(78)
    assign n115 = n6 ? 1'b0 : m_a1[6];   // pipeline_interface.v(78)
    assign n116 = n6 ? 1'b0 : m_a1[5];   // pipeline_interface.v(78)
    assign n117 = n6 ? 1'b0 : m_a1[4];   // pipeline_interface.v(78)
    assign n118 = n6 ? 1'b0 : m_a1[3];   // pipeline_interface.v(78)
    assign n119 = n6 ? 1'b0 : m_a1[2];   // pipeline_interface.v(78)
    assign n120 = n6 ? 1'b0 : m_a1[1];   // pipeline_interface.v(78)
    assign n121 = n6 ? 1'b0 : m_a1[0];   // pipeline_interface.v(78)
    assign n122 = n6 ? 1'b0 : m_a2[31];   // pipeline_interface.v(78)
    assign n123 = n6 ? 1'b0 : m_a2[30];   // pipeline_interface.v(78)
    assign n124 = n6 ? 1'b0 : m_a2[29];   // pipeline_interface.v(78)
    assign n125 = n6 ? 1'b0 : m_a2[28];   // pipeline_interface.v(78)
    assign n126 = n6 ? 1'b0 : m_a2[27];   // pipeline_interface.v(78)
    assign n127 = n6 ? 1'b0 : m_a2[26];   // pipeline_interface.v(78)
    assign n128 = n6 ? 1'b0 : m_a2[25];   // pipeline_interface.v(78)
    assign n129 = n6 ? 1'b0 : m_a2[24];   // pipeline_interface.v(78)
    assign n130 = n6 ? 1'b0 : m_a2[23];   // pipeline_interface.v(78)
    assign n131 = n6 ? 1'b0 : m_a2[22];   // pipeline_interface.v(78)
    assign n132 = n6 ? 1'b0 : m_a2[21];   // pipeline_interface.v(78)
    assign n133 = n6 ? 1'b0 : m_a2[20];   // pipeline_interface.v(78)
    assign n134 = n6 ? 1'b0 : m_a2[19];   // pipeline_interface.v(78)
    assign n135 = n6 ? 1'b0 : m_a2[18];   // pipeline_interface.v(78)
    assign n136 = n6 ? 1'b0 : m_a2[17];   // pipeline_interface.v(78)
    assign n137 = n6 ? 1'b0 : m_a2[16];   // pipeline_interface.v(78)
    assign n138 = n6 ? 1'b0 : m_a2[15];   // pipeline_interface.v(78)
    assign n139 = n6 ? 1'b0 : m_a2[14];   // pipeline_interface.v(78)
    assign n140 = n6 ? 1'b0 : m_a2[13];   // pipeline_interface.v(78)
    assign n141 = n6 ? 1'b0 : m_a2[12];   // pipeline_interface.v(78)
    assign n142 = n6 ? 1'b0 : m_a2[11];   // pipeline_interface.v(78)
    assign n143 = n6 ? 1'b0 : m_a2[10];   // pipeline_interface.v(78)
    assign n144 = n6 ? 1'b0 : m_a2[9];   // pipeline_interface.v(78)
    assign n145 = n6 ? 1'b0 : m_a2[8];   // pipeline_interface.v(78)
    assign n146 = n6 ? 1'b0 : m_a2[7];   // pipeline_interface.v(78)
    assign n147 = n6 ? 1'b0 : m_a2[6];   // pipeline_interface.v(78)
    assign n148 = n6 ? 1'b0 : m_a2[5];   // pipeline_interface.v(78)
    assign n149 = n6 ? 1'b0 : m_a2[4];   // pipeline_interface.v(78)
    assign n150 = n6 ? 1'b0 : m_a2[3];   // pipeline_interface.v(78)
    assign n151 = n6 ? 1'b0 : m_a2[2];   // pipeline_interface.v(78)
    assign n152 = n6 ? 1'b0 : m_a2[1];   // pipeline_interface.v(78)
    assign n153 = n6 ? 1'b0 : m_a2[0];   // pipeline_interface.v(78)
    assign n154 = n6 ? 1'b0 : m_r1_op[3];   // pipeline_interface.v(78)
    assign n155 = n6 ? 1'b0 : m_r1_op[2];   // pipeline_interface.v(78)
    assign n156 = n6 ? 1'b0 : m_r1_op[1];   // pipeline_interface.v(78)
    assign n157 = n6 ? 1'b0 : m_r1_op[0];   // pipeline_interface.v(78)
    assign n158 = n6 ? 1'b0 : m_r2_op[3];   // pipeline_interface.v(78)
    assign n159 = n6 ? 1'b0 : m_r2_op[2];   // pipeline_interface.v(78)
    assign n160 = n6 ? 1'b0 : m_r2_op[1];   // pipeline_interface.v(78)
    assign n161 = n6 ? 1'b0 : m_r2_op[0];   // pipeline_interface.v(78)
    assign n162 = n6 ? 1'b0 : r_a1[4];   // pipeline_interface.v(78)
    assign n163 = n6 ? 1'b0 : r_a1[3];   // pipeline_interface.v(78)
    assign n164 = n6 ? 1'b0 : r_a1[2];   // pipeline_interface.v(78)
    assign n165 = n6 ? 1'b0 : r_a1[1];   // pipeline_interface.v(78)
    assign n166 = n6 ? 1'b0 : r_a1[0];   // pipeline_interface.v(78)
    assign n167 = n6 ? 1'b0 : r_a2[4];   // pipeline_interface.v(78)
    assign n168 = n6 ? 1'b0 : r_a2[3];   // pipeline_interface.v(78)
    assign n169 = n6 ? 1'b0 : r_a2[2];   // pipeline_interface.v(78)
    assign n170 = n6 ? 1'b0 : r_a2[1];   // pipeline_interface.v(78)
    assign n171 = n6 ? 1'b0 : r_a2[0];   // pipeline_interface.v(78)
    assign n172 = n6 ? 1'b0 : r_op[3];   // pipeline_interface.v(78)
    assign n173 = n6 ? 1'b0 : r_op[2];   // pipeline_interface.v(78)
    assign n174 = n6 ? 1'b0 : r_op[1];   // pipeline_interface.v(78)
    assign n175 = n6 ? 1'b0 : r_op[0];   // pipeline_interface.v(78)
    VERIFIC_DFFRS i178 (.d(n9), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[30]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i179 (.d(n10), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[29]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i180 (.d(n11), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[28]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i181 (.d(n12), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[27]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i182 (.d(n13), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[26]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i183 (.d(n14), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[25]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i184 (.d(n15), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[24]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i185 (.d(n16), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[23]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i186 (.d(n17), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[22]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i187 (.d(n18), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[21]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i188 (.d(n19), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[20]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i189 (.d(n20), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[19]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i190 (.d(n21), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[18]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i191 (.d(n22), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[17]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i192 (.d(n23), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[16]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i193 (.d(n24), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[15]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i194 (.d(n25), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[14]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i195 (.d(n26), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[13]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i196 (.d(n27), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[12]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i197 (.d(n28), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[11]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i198 (.d(n29), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[10]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i199 (.d(n30), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[9]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i200 (.d(n31), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[8]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i201 (.d(n32), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[7]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i202 (.d(n33), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[6]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i203 (.d(n34), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[5]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i204 (.d(n35), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[4]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i205 (.d(n36), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[3]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i206 (.d(n37), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[2]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i207 (.d(n38), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[1]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i208 (.d(n39), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[0]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i209 (.d(n40), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[31]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i210 (.d(n41), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[30]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i211 (.d(n42), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[29]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i212 (.d(n43), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[28]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i213 (.d(n44), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[27]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i214 (.d(n45), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[26]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i215 (.d(n46), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[25]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i216 (.d(n47), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[24]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i217 (.d(n48), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[23]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i218 (.d(n49), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[22]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i219 (.d(n50), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[21]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i220 (.d(n51), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[20]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i221 (.d(n52), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[19]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i222 (.d(n53), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[18]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i223 (.d(n54), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[17]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i224 (.d(n55), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[16]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i225 (.d(n56), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[15]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i226 (.d(n57), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[14]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i227 (.d(n58), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[13]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i228 (.d(n59), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[12]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i229 (.d(n60), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[11]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i230 (.d(n61), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[10]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i231 (.d(n62), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[9]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i232 (.d(n63), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[8]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i233 (.d(n64), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[7]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i234 (.d(n65), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[6]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i235 (.d(n66), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[5]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i236 (.d(n67), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[4]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i237 (.d(n68), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[3]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i238 (.d(n69), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[2]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i239 (.d(n70), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[1]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i240 (.d(n71), .clk(clk), .s(1'b0), .r(rst), .q(qe_b[0]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i241 (.d(n72), .clk(clk), .s(1'b0), .r(rst), .q(qe_alu_op[7]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i242 (.d(n73), .clk(clk), .s(1'b0), .r(rst), .q(qe_alu_op[6]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i243 (.d(n74), .clk(clk), .s(1'b0), .r(rst), .q(qe_alu_op[5]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i244 (.d(n75), .clk(clk), .s(1'b0), .r(rst), .q(qe_alu_op[4]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i245 (.d(n76), .clk(clk), .s(1'b0), .r(rst), .q(qe_alu_op[3]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i246 (.d(n77), .clk(clk), .s(1'b0), .r(rst), .q(qe_alu_op[2]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i247 (.d(n78), .clk(clk), .s(1'b0), .r(rst), .q(qe_alu_op[1]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i248 (.d(n79), .clk(clk), .s(1'b0), .r(rst), .q(qe_alu_op[0]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i249 (.d(n80), .clk(clk), .s(1'b0), .r(rst), .q(qe_cond[3]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i250 (.d(n81), .clk(clk), .s(1'b0), .r(rst), .q(qe_cond[2]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i251 (.d(n82), .clk(clk), .s(1'b0), .r(rst), .q(qe_cond[1]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i252 (.d(n83), .clk(clk), .s(1'b0), .r(rst), .q(qe_cond[0]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i253 (.d(n84), .clk(clk), .s(1'b0), .r(rst), .q(qe_write_flags[3]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i254 (.d(n85), .clk(clk), .s(1'b0), .r(rst), .q(qe_write_flags[2]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i255 (.d(n86), .clk(clk), .s(1'b0), .r(rst), .q(qe_write_flags[1]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i256 (.d(n87), .clk(clk), .s(1'b0), .r(rst), .q(qe_write_flags[0]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i257 (.d(n88), .clk(clk), .s(1'b0), .r(rst), .q(qe_swp));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i258 (.d(n89), .clk(clk), .s(1'b0), .r(rst), .q(qe_is_cond));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i259 (.d(n90), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[31]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i260 (.d(n91), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[30]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i261 (.d(n92), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[29]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i262 (.d(n93), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[28]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i263 (.d(n94), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[27]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i264 (.d(n95), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[26]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i265 (.d(n96), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[25]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i266 (.d(n97), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[24]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i267 (.d(n98), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[23]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i268 (.d(n99), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[22]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i269 (.d(n100), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[21]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i270 (.d(n101), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[20]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i271 (.d(n102), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[19]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i272 (.d(n103), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[18]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i273 (.d(n104), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[17]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i274 (.d(n105), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[16]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i275 (.d(n106), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[15]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i276 (.d(n107), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[14]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i277 (.d(n108), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[13]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i278 (.d(n109), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[12]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i279 (.d(n110), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[11]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i280 (.d(n111), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[10]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i281 (.d(n112), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[9]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i282 (.d(n113), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[8]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i283 (.d(n114), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[7]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i284 (.d(n115), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[6]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i285 (.d(n116), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[5]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i286 (.d(n117), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[4]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i287 (.d(n118), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[3]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i288 (.d(n119), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[2]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i289 (.d(n120), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[1]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i290 (.d(n121), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[0]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i291 (.d(n122), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[31]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i292 (.d(n123), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[30]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i293 (.d(n124), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[29]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i294 (.d(n125), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[28]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i295 (.d(n126), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[27]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i296 (.d(n127), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[26]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i297 (.d(n128), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[25]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i298 (.d(n129), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[24]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i299 (.d(n130), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[23]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i300 (.d(n131), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[22]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i301 (.d(n132), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[21]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i302 (.d(n133), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[20]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i303 (.d(n134), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[19]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i304 (.d(n135), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[18]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i305 (.d(n136), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[17]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i306 (.d(n137), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[16]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i307 (.d(n138), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[15]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i308 (.d(n139), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[14]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i309 (.d(n140), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[13]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i310 (.d(n141), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[12]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i311 (.d(n142), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[11]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i312 (.d(n143), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[10]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i313 (.d(n144), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[9]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i314 (.d(n145), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[8]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i315 (.d(n146), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[7]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i316 (.d(n147), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[6]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i317 (.d(n148), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[5]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i318 (.d(n149), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[4]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i319 (.d(n150), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[3]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i320 (.d(n151), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[2]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i321 (.d(n152), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[1]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i322 (.d(n153), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[0]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i323 (.d(n154), .clk(clk), .s(1'b0), .r(rst), .q(qm_r1_op[3]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i324 (.d(n155), .clk(clk), .s(1'b0), .r(rst), .q(qm_r1_op[2]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i325 (.d(n156), .clk(clk), .s(1'b0), .r(rst), .q(qm_r1_op[1]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i326 (.d(n157), .clk(clk), .s(1'b0), .r(rst), .q(qm_r1_op[0]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i327 (.d(n158), .clk(clk), .s(1'b0), .r(rst), .q(qm_r2_op[3]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i328 (.d(n159), .clk(clk), .s(1'b0), .r(rst), .q(qm_r2_op[2]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i329 (.d(n160), .clk(clk), .s(1'b0), .r(rst), .q(qm_r2_op[1]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i330 (.d(n161), .clk(clk), .s(1'b0), .r(rst), .q(qm_r2_op[0]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i331 (.d(n162), .clk(clk), .s(1'b0), .r(rst), .q(qr_a1[4]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i332 (.d(n163), .clk(clk), .s(1'b0), .r(rst), .q(qr_a1[3]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i333 (.d(n164), .clk(clk), .s(1'b0), .r(rst), .q(qr_a1[2]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i334 (.d(n165), .clk(clk), .s(1'b0), .r(rst), .q(qr_a1[1]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i335 (.d(n166), .clk(clk), .s(1'b0), .r(rst), .q(qr_a1[0]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i336 (.d(n167), .clk(clk), .s(1'b0), .r(rst), .q(qr_a2[4]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i337 (.d(n168), .clk(clk), .s(1'b0), .r(rst), .q(qr_a2[3]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i338 (.d(n169), .clk(clk), .s(1'b0), .r(rst), .q(qr_a2[2]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i339 (.d(n170), .clk(clk), .s(1'b0), .r(rst), .q(qr_a2[1]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i340 (.d(n171), .clk(clk), .s(1'b0), .r(rst), .q(qr_a2[0]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i341 (.d(n172), .clk(clk), .s(1'b0), .r(rst), .q(qr_op[3]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i342 (.d(n173), .clk(clk), .s(1'b0), .r(rst), .q(qr_op[2]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i343 (.d(n174), .clk(clk), .s(1'b0), .r(rst), .q(qr_op[1]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i344 (.d(n175), .clk(clk), .s(1'b0), .r(rst), .q(qr_op[0]));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i346 (.d(d_pcincr), .clk(clk), .s(rst), .r(1'b0), 
            .q(qd_pcincr));   // pipeline_interface.v(60)
    VERIFIC_DFFRS i177 (.d(n8), .clk(clk), .s(1'b0), .r(rst), .q(qe_a[31]));   // pipeline_interface.v(60)
    
endmodule

//
// Verific Verilog Description of module execute
//

module execute (r1, r2, cres, n, z, c, v, cc, a, b, alu_op, 
            is_cond, cond, write_flags, st, swp, clk, rst);   // execute.v(78)
    output [31:0]r1;   // execute.v(88)
    output [31:0]r2;   // execute.v(88)
    output cres;   // execute.v(91)
    output n;   // execute.v(89)
    output z;   // execute.v(89)
    output c;   // execute.v(89)
    output v;   // execute.v(89)
    output cc;   // execute.v(90)
    input [31:0]a;   // execute.v(79)
    input [31:0]b;   // execute.v(79)
    input [7:0]alu_op;   // execute.v(81)
    input is_cond;   // execute.v(82)
    input [3:0]cond;   // execute.v(83)
    input [3:0]write_flags;   // execute.v(84)
    input [31:0]st;   // execute.v(80)
    input swp;   // execute.v(85)
    input clk;   // execute.v(86)
    input rst;   // execute.v(86)
    
    wire [31:0]ra;   // execute.v(93)
    wire [31:0]rb;   // execute.v(94)
    wire [31:0]alu_q1;   // execute.v(96)
    wire [31:0]alu_q2;   // execute.v(96)
    wire alu_n;   // execute.v(97)
    wire alu_z;   // execute.v(97)
    wire alu_c;   // execute.v(97)
    wire alu_v;   // execute.v(97)
    wire cond_res;   // execute.v(102)
    
    wire n137, n138, n145;
    
    assign ra[31] = swp ? b[31] : a[31];   // execute.v(93)
    assign ra[30] = swp ? b[30] : a[30];   // execute.v(93)
    assign ra[29] = swp ? b[29] : a[29];   // execute.v(93)
    assign ra[28] = swp ? b[28] : a[28];   // execute.v(93)
    assign ra[27] = swp ? b[27] : a[27];   // execute.v(93)
    assign ra[26] = swp ? b[26] : a[26];   // execute.v(93)
    assign ra[25] = swp ? b[25] : a[25];   // execute.v(93)
    assign ra[24] = swp ? b[24] : a[24];   // execute.v(93)
    assign ra[23] = swp ? b[23] : a[23];   // execute.v(93)
    assign ra[22] = swp ? b[22] : a[22];   // execute.v(93)
    assign ra[21] = swp ? b[21] : a[21];   // execute.v(93)
    assign ra[20] = swp ? b[20] : a[20];   // execute.v(93)
    assign ra[19] = swp ? b[19] : a[19];   // execute.v(93)
    assign ra[18] = swp ? b[18] : a[18];   // execute.v(93)
    assign ra[17] = swp ? b[17] : a[17];   // execute.v(93)
    assign ra[16] = swp ? b[16] : a[16];   // execute.v(93)
    assign ra[15] = swp ? b[15] : a[15];   // execute.v(93)
    assign ra[14] = swp ? b[14] : a[14];   // execute.v(93)
    assign ra[13] = swp ? b[13] : a[13];   // execute.v(93)
    assign ra[12] = swp ? b[12] : a[12];   // execute.v(93)
    assign ra[11] = swp ? b[11] : a[11];   // execute.v(93)
    assign ra[10] = swp ? b[10] : a[10];   // execute.v(93)
    assign ra[9] = swp ? b[9] : a[9];   // execute.v(93)
    assign ra[8] = swp ? b[8] : a[8];   // execute.v(93)
    assign ra[7] = swp ? b[7] : a[7];   // execute.v(93)
    assign ra[6] = swp ? b[6] : a[6];   // execute.v(93)
    assign ra[5] = swp ? b[5] : a[5];   // execute.v(93)
    assign ra[4] = swp ? b[4] : a[4];   // execute.v(93)
    assign ra[3] = swp ? b[3] : a[3];   // execute.v(93)
    assign ra[2] = swp ? b[2] : a[2];   // execute.v(93)
    assign ra[1] = swp ? b[1] : a[1];   // execute.v(93)
    assign ra[0] = swp ? b[0] : a[0];   // execute.v(93)
    assign rb[31] = swp ? a[31] : b[31];   // execute.v(94)
    assign rb[30] = swp ? a[30] : b[30];   // execute.v(94)
    assign rb[29] = swp ? a[29] : b[29];   // execute.v(94)
    assign rb[28] = swp ? a[28] : b[28];   // execute.v(94)
    assign rb[27] = swp ? a[27] : b[27];   // execute.v(94)
    assign rb[26] = swp ? a[26] : b[26];   // execute.v(94)
    assign rb[25] = swp ? a[25] : b[25];   // execute.v(94)
    assign rb[24] = swp ? a[24] : b[24];   // execute.v(94)
    assign rb[23] = swp ? a[23] : b[23];   // execute.v(94)
    assign rb[22] = swp ? a[22] : b[22];   // execute.v(94)
    assign rb[21] = swp ? a[21] : b[21];   // execute.v(94)
    assign rb[20] = swp ? a[20] : b[20];   // execute.v(94)
    assign rb[19] = swp ? a[19] : b[19];   // execute.v(94)
    assign rb[18] = swp ? a[18] : b[18];   // execute.v(94)
    assign rb[17] = swp ? a[17] : b[17];   // execute.v(94)
    assign rb[16] = swp ? a[16] : b[16];   // execute.v(94)
    assign rb[15] = swp ? a[15] : b[15];   // execute.v(94)
    assign rb[14] = swp ? a[14] : b[14];   // execute.v(94)
    assign rb[13] = swp ? a[13] : b[13];   // execute.v(94)
    assign rb[12] = swp ? a[12] : b[12];   // execute.v(94)
    assign rb[11] = swp ? a[11] : b[11];   // execute.v(94)
    assign rb[10] = swp ? a[10] : b[10];   // execute.v(94)
    assign rb[9] = swp ? a[9] : b[9];   // execute.v(94)
    assign rb[8] = swp ? a[8] : b[8];   // execute.v(94)
    assign rb[7] = swp ? a[7] : b[7];   // execute.v(94)
    assign rb[6] = swp ? a[6] : b[6];   // execute.v(94)
    assign rb[5] = swp ? a[5] : b[5];   // execute.v(94)
    assign rb[4] = swp ? a[4] : b[4];   // execute.v(94)
    assign rb[3] = swp ? a[3] : b[3];   // execute.v(94)
    assign rb[2] = swp ? a[2] : b[2];   // execute.v(94)
    assign rb[1] = swp ? a[1] : b[1];   // execute.v(94)
    assign rb[0] = swp ? a[0] : b[0];   // execute.v(94)
    alu32_2x2 alu0 (.q0({alu_q1}), .q1({alu_q2}), .st({alu_n, alu_z, 
            alu_c, alu_v}), .a({ra}), .b({rb}), .op({alu_op}));   // execute.v(99)
    cond_calc cond0 (.cr(cond_res), .cc({cond}), .n(st[3]), .z(st[2]), 
            .c(st[1]), .v(st[0]));   // execute.v(103)
    or (n137, write_flags[3], write_flags[2], write_flags[1], write_flags[0]) ;   // execute.v(105)
    and (n138, is_cond, cond_res) ;   // execute.v(105)
    and (cc, n137, n138) ;   // execute.v(105)
    assign n = write_flags[3] ? alu_n : st[3];   // execute.v(106)
    assign z = write_flags[2] ? alu_z : st[2];   // execute.v(107)
    assign c = write_flags[1] ? alu_c : st[1];   // execute.v(108)
    assign v = write_flags[0] ? alu_v : st[0];   // execute.v(109)
    assign n145 = is_cond ? cond_res : 1'b1;   // execute.v(121)
    VERIFIC_DFFRS i78 (.d(alu_q1[30]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[30]));   // execute.v(117)
    VERIFIC_DFFRS i79 (.d(alu_q1[29]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[29]));   // execute.v(117)
    VERIFIC_DFFRS i80 (.d(alu_q1[28]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[28]));   // execute.v(117)
    VERIFIC_DFFRS i81 (.d(alu_q1[27]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[27]));   // execute.v(117)
    VERIFIC_DFFRS i82 (.d(alu_q1[26]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[26]));   // execute.v(117)
    VERIFIC_DFFRS i83 (.d(alu_q1[25]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[25]));   // execute.v(117)
    VERIFIC_DFFRS i84 (.d(alu_q1[24]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[24]));   // execute.v(117)
    VERIFIC_DFFRS i85 (.d(alu_q1[23]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[23]));   // execute.v(117)
    VERIFIC_DFFRS i86 (.d(alu_q1[22]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[22]));   // execute.v(117)
    VERIFIC_DFFRS i87 (.d(alu_q1[21]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[21]));   // execute.v(117)
    VERIFIC_DFFRS i88 (.d(alu_q1[20]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[20]));   // execute.v(117)
    VERIFIC_DFFRS i89 (.d(alu_q1[19]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[19]));   // execute.v(117)
    VERIFIC_DFFRS i90 (.d(alu_q1[18]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[18]));   // execute.v(117)
    VERIFIC_DFFRS i91 (.d(alu_q1[17]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[17]));   // execute.v(117)
    VERIFIC_DFFRS i92 (.d(alu_q1[16]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[16]));   // execute.v(117)
    VERIFIC_DFFRS i93 (.d(alu_q1[15]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[15]));   // execute.v(117)
    VERIFIC_DFFRS i94 (.d(alu_q1[14]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[14]));   // execute.v(117)
    VERIFIC_DFFRS i95 (.d(alu_q1[13]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[13]));   // execute.v(117)
    VERIFIC_DFFRS i96 (.d(alu_q1[12]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[12]));   // execute.v(117)
    VERIFIC_DFFRS i97 (.d(alu_q1[11]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[11]));   // execute.v(117)
    VERIFIC_DFFRS i98 (.d(alu_q1[10]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[10]));   // execute.v(117)
    VERIFIC_DFFRS i99 (.d(alu_q1[9]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[9]));   // execute.v(117)
    VERIFIC_DFFRS i100 (.d(alu_q1[8]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[8]));   // execute.v(117)
    VERIFIC_DFFRS i101 (.d(alu_q1[7]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[7]));   // execute.v(117)
    VERIFIC_DFFRS i102 (.d(alu_q1[6]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[6]));   // execute.v(117)
    VERIFIC_DFFRS i103 (.d(alu_q1[5]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[5]));   // execute.v(117)
    VERIFIC_DFFRS i104 (.d(alu_q1[4]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[4]));   // execute.v(117)
    VERIFIC_DFFRS i105 (.d(alu_q1[3]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[3]));   // execute.v(117)
    VERIFIC_DFFRS i106 (.d(alu_q1[2]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[2]));   // execute.v(117)
    VERIFIC_DFFRS i107 (.d(alu_q1[1]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[1]));   // execute.v(117)
    VERIFIC_DFFRS i108 (.d(alu_q1[0]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[0]));   // execute.v(117)
    VERIFIC_DFFRS i109 (.d(alu_q2[31]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[31]));   // execute.v(117)
    VERIFIC_DFFRS i110 (.d(alu_q2[30]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[30]));   // execute.v(117)
    VERIFIC_DFFRS i111 (.d(alu_q2[29]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[29]));   // execute.v(117)
    VERIFIC_DFFRS i112 (.d(alu_q2[28]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[28]));   // execute.v(117)
    VERIFIC_DFFRS i113 (.d(alu_q2[27]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[27]));   // execute.v(117)
    VERIFIC_DFFRS i114 (.d(alu_q2[26]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[26]));   // execute.v(117)
    VERIFIC_DFFRS i115 (.d(alu_q2[25]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[25]));   // execute.v(117)
    VERIFIC_DFFRS i116 (.d(alu_q2[24]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[24]));   // execute.v(117)
    VERIFIC_DFFRS i117 (.d(alu_q2[23]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[23]));   // execute.v(117)
    VERIFIC_DFFRS i118 (.d(alu_q2[22]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[22]));   // execute.v(117)
    VERIFIC_DFFRS i119 (.d(alu_q2[21]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[21]));   // execute.v(117)
    VERIFIC_DFFRS i120 (.d(alu_q2[20]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[20]));   // execute.v(117)
    VERIFIC_DFFRS i121 (.d(alu_q2[19]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[19]));   // execute.v(117)
    VERIFIC_DFFRS i122 (.d(alu_q2[18]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[18]));   // execute.v(117)
    VERIFIC_DFFRS i123 (.d(alu_q2[17]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[17]));   // execute.v(117)
    VERIFIC_DFFRS i124 (.d(alu_q2[16]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[16]));   // execute.v(117)
    VERIFIC_DFFRS i125 (.d(alu_q2[15]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[15]));   // execute.v(117)
    VERIFIC_DFFRS i126 (.d(alu_q2[14]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[14]));   // execute.v(117)
    VERIFIC_DFFRS i127 (.d(alu_q2[13]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[13]));   // execute.v(117)
    VERIFIC_DFFRS i128 (.d(alu_q2[12]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[12]));   // execute.v(117)
    VERIFIC_DFFRS i129 (.d(alu_q2[11]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[11]));   // execute.v(117)
    VERIFIC_DFFRS i130 (.d(alu_q2[10]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[10]));   // execute.v(117)
    VERIFIC_DFFRS i131 (.d(alu_q2[9]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[9]));   // execute.v(117)
    VERIFIC_DFFRS i132 (.d(alu_q2[8]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[8]));   // execute.v(117)
    VERIFIC_DFFRS i133 (.d(alu_q2[7]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[7]));   // execute.v(117)
    VERIFIC_DFFRS i134 (.d(alu_q2[6]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[6]));   // execute.v(117)
    VERIFIC_DFFRS i135 (.d(alu_q2[5]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[5]));   // execute.v(117)
    VERIFIC_DFFRS i136 (.d(alu_q2[4]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[4]));   // execute.v(117)
    VERIFIC_DFFRS i137 (.d(alu_q2[3]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[3]));   // execute.v(117)
    VERIFIC_DFFRS i138 (.d(alu_q2[2]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[2]));   // execute.v(117)
    VERIFIC_DFFRS i139 (.d(alu_q2[1]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[1]));   // execute.v(117)
    VERIFIC_DFFRS i140 (.d(alu_q2[0]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r2[0]));   // execute.v(117)
    VERIFIC_DFFRS i141 (.d(n145), .clk(clk), .s(1'b0), .r(rst), .q(cres));   // execute.v(117)
    VERIFIC_DFFRS i77 (.d(alu_q1[31]), .clk(clk), .s(1'b0), .r(rst), 
            .q(r1[31]));   // execute.v(117)
    
endmodule

//
// Verific Verilog Description of module alu32_2x2
//

module alu32_2x2 (q0, q1, st, a, b, op);   // alu.v(62)
    output [31:0]q0;   // alu.v(64)
    output [31:0]q1;   // alu.v(64)
    output [3:0]st;   // alu.v(68)
    input [31:0]a;   // alu.v(63)
    input [31:0]b;   // alu.v(63)
    input [7:0]op;   // alu.v(67)
    
    wire [31:0]addsub;   // alu.v(70)
    wire [31:0]addsub_a;   // alu.v(71)
    wire [31:0]addsub_b;   // alu.v(71)
    wire subtract;   // alu.v(73)
    wire [3:0]addsub_st;   // alu.v(75)
    wire [31:0]shift;   // alu.v(78)
    wire rotate;   // alu.v(80)
    wire left;   // alu.v(80)
    wire arithmetic;   // alu.v(80)
    wire [3:0]shift_st;   // alu.v(82)
    wire [31:0]mull;   // alu.v(84)
    wire [31:0]mulh;   // alu.v(84)
    wire [3:0]mul_st;   // alu.v(87)
    wire [31:0]bws;   // alu.v(89)
    wire [2:0]b_op;   // alu.v(91)
    wire [3:0]bws_st;   // alu.v(93)
    
    wire n172, n173, n174, n175, n176, n179, n180, n181, n184, 
        n187, n191, n192, n193, n196, n199, n203, n206, n210, 
        n214, n219, n220, n221, n224, n225, n226, n227, n228, 
        n354, n434, n435, n438, n629, n630, n631, n634, n635, 
        n638, n639, n641, n642, n643, n646, n647, n650, n651, 
        n655, n657, n661, n667, n673, n679, n685, n691, n697, 
        n703, n709, n715, n721, n727, n733, n739, n745, n751, 
        n757, n763, n769, n775, n781, n787, n793, n799, n805, 
        n811, n817, n823, n829, n835, n841, n847, n849, n853, 
        n859, n865, n871, n877, n883, n889, n895, n901, n907, 
        n913, n919, n925, n931, n937, n943, n949, n955, n961, 
        n967, n973, n979, n985, n991, n997, n1003, n1009, n1015, 
        n1021, n1027, n1033, n1039, n1045, n1051, n1057, n1063, 
        n1065, n1069, n1071, n1075, n1081, n1087, n1093, n1099, 
        n1105, n1111, n1117, n1123, n1129, n1135, n1141, n1147, 
        n1153, n1159, n1165, n1171, n1177, n1183, n1189, n1195, 
        n1201, n1207, n1213, n1219, n1225, n1231, n1237, n1243, 
        n1249, n1255, n1261, n1267, n1273, n1279, n1285, n1291, 
        n1297, n1303, n1309, n1315, n1321, n1327, n1333, n1339, 
        n1345, n1351, n1357, n1363, n1369, n1375, n1381, n1387, 
        n1393, n1399, n1405, n1411, n1417, n1423, n1429, n1435, 
        n1441, n1447, n1453, n1455, n1459, n1461, n1465, n1467, 
        n1471, n1473, n1477, n1479, n1483, n1485;
    
    addsub_32 as0 (.q({addsub}), .a({addsub_a}), .b({addsub_b}), .sub(subtract), 
            .ov(addsub_st[1]), .sov(addsub_st[0]), .z(addsub_st[2]));   // alu.v(74)
    bshift_32 sh0 (.q({shift}), .ov(shift_st[1]), .z(shift_st[2]), .a({a}), 
            .b({b[4:0]}), .rotate(rotate), .left(left), .arith(arithmetic));   // alu.v(81)
    mul_32 mul0 (.q1({mull}), .q2({mulh}), .ov(mul_st[1]), .z(mul_st[2]), 
           .a({a}), .b({b}));   // alu.v(86)
    bitwise_32 bw0 (.q({bws}), .z(bws_st[2]), .a({a}), .b({b}), .op({b_op}));   // alu.v(92)
    nor (n172, op[7], op[6], op[5], op[4], op[3], op[2], op[1], 
            op[0]) ;   // alu.v(98)
    not (n173, op[0]) ;   // alu.v(104)
    nor (n174, op[7], op[6], op[5], op[4], op[3], op[2], op[1], 
        n173) ;   // alu.v(104)
    not (n175, op[1]) ;   // alu.v(113)
    nor (n176, op[7], op[6], op[5], op[4], op[3], op[2], n175, 
        op[0]) ;   // alu.v(113)
    nor (n179, op[7], op[6], op[5], op[4], op[3], op[2], n175, 
        n173) ;   // alu.v(122)
    not (n180, op[2]) ;   // alu.v(131)
    nor (n181, op[7], op[6], op[5], op[4], op[3], n180, op[1], 
        op[0]) ;   // alu.v(131)
    nor (n184, op[7], op[6], op[5], op[4], op[3], n180, op[1], 
        n173) ;   // alu.v(137)
    nor (n187, op[7], op[6], op[5], op[4], op[3], n180, n175, 
        op[0]) ;   // alu.v(146)
    nor (n191, op[7], op[6], op[5], op[4], op[3], n180, n175, 
        n173) ;   // alu.v(155)
    not (n192, op[3]) ;   // alu.v(164)
    nor (n193, op[7], op[6], op[5], op[4], n192, op[2], op[1], 
        op[0]) ;   // alu.v(164)
    nor (n196, op[7], op[6], op[5], op[4], n192, op[2], op[1], 
        n173) ;   // alu.v(173)
    nor (n199, op[7], op[6], op[5], op[4], n192, op[2], n175, 
        op[0]) ;   // alu.v(182)
    nor (n203, op[7], op[6], op[5], op[4], n192, op[2], n175, 
        n173) ;   // alu.v(191)
    nor (n206, op[7], op[6], op[5], op[4], n192, n180, op[1], 
        op[0]) ;   // alu.v(198)
    nor (n210, op[7], op[6], op[5], op[4], n192, n180, op[1], 
        n173) ;   // alu.v(205)
    nor (n214, op[7], op[6], op[5], op[4], n192, n180, n175, 
        op[0]) ;   // alu.v(212)
    nor (n219, op[7], op[6], op[5], op[4], n192, n180, n175, 
        n173) ;   // alu.v(219)
    not (n220, op[4]) ;   // alu.v(226)
    nor (n221, op[7], op[6], op[5], n220, op[3], op[2], op[1], 
        op[0]) ;   // alu.v(226)
    nor (n224, op[7], op[6], op[5], n220, op[3], op[2], op[1], 
        n173) ;   // alu.v(233)
    nor (n225, n172, n174, n176, n179, n181, n184, n187, n191, 
        n193, n196, n199, n203, n206, n210, n214, n219, n221, 
        n224) ;   // alu.v(97)
    or (n226, n174, n176, n179) ;   // alu.v(97)
    or (n227, n184, n187, n191, n193, n196, n199) ;   // alu.v(97)
    or (n228, n203, n206, n210, n214, n219, n221, n224) ;   // alu.v(97)
    or (n354, n174, n176, n179, n184, n187, n191, n193, n196, 
        n199, n203, n206, n210, n214, n219, n221, n224) ;   // alu.v(97)
    or (n434, n172, n181, n184, n187, n191, n193, n196, n199, 
        n203, n206, n210, n214, n219, n221, n224, n225) ;   // alu.v(97)
    or (n435, n176, n179) ;   // alu.v(97)
    or (n438, n174, n176) ;   // alu.v(97)
    or (n629, n172, n174, n176, n179, n181, n203, n206, n210, 
        n214, n219, n221, n224, n225) ;   // alu.v(97)
    or (n630, n184, n187, n191, n193) ;   // alu.v(97)
    or (n631, n196, n199) ;   // alu.v(97)
    or (n634, n184, n191, n196) ;   // alu.v(97)
    or (n635, n187, n193, n199) ;   // alu.v(97)
    or (n638, n184, n187, n196, n199) ;   // alu.v(97)
    or (n639, n191, n193) ;   // alu.v(97)
    or (n641, n172, n174, n176, n179, n181, n184, n187, n191, 
        n193, n196, n199, n225) ;   // alu.v(97)
    or (n642, n203, n206, n210, n214) ;   // alu.v(97)
    or (n643, n219, n221, n224) ;   // alu.v(97)
    or (n646, n203, n206, n219, n221) ;   // alu.v(97)
    or (n647, n210, n214, n224) ;   // alu.v(97)
    or (n650, n203, n210, n219, n224) ;   // alu.v(97)
    or (n651, n206, n214, n221) ;   // alu.v(97)
    Select_6 Select_486 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[31], addsub[31], mull[31], shift[31], bws[31], 
            1'bx}), .o(n655));   // alu.v(97)
    Select_6 Select_488 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({6'b111110}), .o(n657));   // alu.v(97)
    assign q0[31] = n657 ? n655 : 1'bz;   // alu.v(96)
    Select_6 Select_492 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[30], addsub[30], mull[30], shift[30], bws[30], 
            1'bx}), .o(n661));   // alu.v(97)
    assign q0[30] = n657 ? n661 : 1'bz;   // alu.v(96)
    Select_6 Select_498 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[29], addsub[29], mull[29], shift[29], bws[29], 
            1'bx}), .o(n667));   // alu.v(97)
    assign q0[29] = n657 ? n667 : 1'bz;   // alu.v(96)
    Select_6 Select_504 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[28], addsub[28], mull[28], shift[28], bws[28], 
            1'bx}), .o(n673));   // alu.v(97)
    assign q0[28] = n657 ? n673 : 1'bz;   // alu.v(96)
    Select_6 Select_510 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[27], addsub[27], mull[27], shift[27], bws[27], 
            1'bx}), .o(n679));   // alu.v(97)
    assign q0[27] = n657 ? n679 : 1'bz;   // alu.v(96)
    Select_6 Select_516 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[26], addsub[26], mull[26], shift[26], bws[26], 
            1'bx}), .o(n685));   // alu.v(97)
    assign q0[26] = n657 ? n685 : 1'bz;   // alu.v(96)
    Select_6 Select_522 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[25], addsub[25], mull[25], shift[25], bws[25], 
            1'bx}), .o(n691));   // alu.v(97)
    assign q0[25] = n657 ? n691 : 1'bz;   // alu.v(96)
    Select_6 Select_528 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[24], addsub[24], mull[24], shift[24], bws[24], 
            1'bx}), .o(n697));   // alu.v(97)
    assign q0[24] = n657 ? n697 : 1'bz;   // alu.v(96)
    Select_6 Select_534 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[23], addsub[23], mull[23], shift[23], bws[23], 
            1'bx}), .o(n703));   // alu.v(97)
    assign q0[23] = n657 ? n703 : 1'bz;   // alu.v(96)
    Select_6 Select_540 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[22], addsub[22], mull[22], shift[22], bws[22], 
            1'bx}), .o(n709));   // alu.v(97)
    assign q0[22] = n657 ? n709 : 1'bz;   // alu.v(96)
    Select_6 Select_546 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[21], addsub[21], mull[21], shift[21], bws[21], 
            1'bx}), .o(n715));   // alu.v(97)
    assign q0[21] = n657 ? n715 : 1'bz;   // alu.v(96)
    Select_6 Select_552 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[20], addsub[20], mull[20], shift[20], bws[20], 
            1'bx}), .o(n721));   // alu.v(97)
    assign q0[20] = n657 ? n721 : 1'bz;   // alu.v(96)
    Select_6 Select_558 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[19], addsub[19], mull[19], shift[19], bws[19], 
            1'bx}), .o(n727));   // alu.v(97)
    assign q0[19] = n657 ? n727 : 1'bz;   // alu.v(96)
    Select_6 Select_564 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[18], addsub[18], mull[18], shift[18], bws[18], 
            1'bx}), .o(n733));   // alu.v(97)
    assign q0[18] = n657 ? n733 : 1'bz;   // alu.v(96)
    Select_6 Select_570 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[17], addsub[17], mull[17], shift[17], bws[17], 
            1'bx}), .o(n739));   // alu.v(97)
    assign q0[17] = n657 ? n739 : 1'bz;   // alu.v(96)
    Select_6 Select_576 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[16], addsub[16], mull[16], shift[16], bws[16], 
            1'bx}), .o(n745));   // alu.v(97)
    assign q0[16] = n657 ? n745 : 1'bz;   // alu.v(96)
    Select_6 Select_582 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[15], addsub[15], mull[15], shift[15], bws[15], 
            1'bx}), .o(n751));   // alu.v(97)
    assign q0[15] = n657 ? n751 : 1'bz;   // alu.v(96)
    Select_6 Select_588 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[14], addsub[14], mull[14], shift[14], bws[14], 
            1'bx}), .o(n757));   // alu.v(97)
    assign q0[14] = n657 ? n757 : 1'bz;   // alu.v(96)
    Select_6 Select_594 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[13], addsub[13], mull[13], shift[13], bws[13], 
            1'bx}), .o(n763));   // alu.v(97)
    assign q0[13] = n657 ? n763 : 1'bz;   // alu.v(96)
    Select_6 Select_600 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[12], addsub[12], mull[12], shift[12], bws[12], 
            1'bx}), .o(n769));   // alu.v(97)
    assign q0[12] = n657 ? n769 : 1'bz;   // alu.v(96)
    Select_6 Select_606 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[11], addsub[11], mull[11], shift[11], bws[11], 
            1'bx}), .o(n775));   // alu.v(97)
    assign q0[11] = n657 ? n775 : 1'bz;   // alu.v(96)
    Select_6 Select_612 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[10], addsub[10], mull[10], shift[10], bws[10], 
            1'bx}), .o(n781));   // alu.v(97)
    assign q0[10] = n657 ? n781 : 1'bz;   // alu.v(96)
    Select_6 Select_618 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[9], addsub[9], mull[9], shift[9], bws[9], 1'bx}), 
            .o(n787));   // alu.v(97)
    assign q0[9] = n657 ? n787 : 1'bz;   // alu.v(96)
    Select_6 Select_624 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[8], addsub[8], mull[8], shift[8], bws[8], 1'bx}), 
            .o(n793));   // alu.v(97)
    assign q0[8] = n657 ? n793 : 1'bz;   // alu.v(96)
    Select_6 Select_630 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[7], addsub[7], mull[7], shift[7], bws[7], 1'bx}), 
            .o(n799));   // alu.v(97)
    assign q0[7] = n657 ? n799 : 1'bz;   // alu.v(96)
    Select_6 Select_636 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[6], addsub[6], mull[6], shift[6], bws[6], 1'bx}), 
            .o(n805));   // alu.v(97)
    assign q0[6] = n657 ? n805 : 1'bz;   // alu.v(96)
    Select_6 Select_642 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[5], addsub[5], mull[5], shift[5], bws[5], 1'bx}), 
            .o(n811));   // alu.v(97)
    assign q0[5] = n657 ? n811 : 1'bz;   // alu.v(96)
    Select_6 Select_648 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[4], addsub[4], mull[4], shift[4], bws[4], 1'bx}), 
            .o(n817));   // alu.v(97)
    assign q0[4] = n657 ? n817 : 1'bz;   // alu.v(96)
    Select_6 Select_654 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[3], addsub[3], mull[3], shift[3], bws[3], 1'bx}), 
            .o(n823));   // alu.v(97)
    assign q0[3] = n657 ? n823 : 1'bz;   // alu.v(96)
    Select_6 Select_660 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[2], addsub[2], mull[2], shift[2], bws[2], 1'bx}), 
            .o(n829));   // alu.v(97)
    assign q0[2] = n657 ? n829 : 1'bz;   // alu.v(96)
    Select_6 Select_666 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[1], addsub[1], mull[1], shift[1], bws[1], 1'bx}), 
            .o(n835));   // alu.v(97)
    assign q0[1] = n657 ? n835 : 1'bz;   // alu.v(96)
    Select_6 Select_672 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({a[0], addsub[0], mull[0], shift[0], bws[0], 1'bx}), 
            .o(n841));   // alu.v(97)
    assign q0[0] = n657 ? n841 : 1'bz;   // alu.v(96)
    Select_4 Select_678 (.sel({n172, n354, n181, n225}), .data({b[31], 
            1'b0, mulh[31], 1'bx}), .o(n847));   // alu.v(97)
    Select_4 Select_680 (.sel({n172, n354, n181, n225}), .data({4'b1110}), 
            .o(n849));   // alu.v(97)
    assign q1[31] = n849 ? n847 : 1'bz;   // alu.v(96)
    Select_4 Select_684 (.sel({n172, n354, n181, n225}), .data({b[30], 
            1'b0, mulh[30], 1'bx}), .o(n853));   // alu.v(97)
    assign q1[30] = n849 ? n853 : 1'bz;   // alu.v(96)
    Select_4 Select_690 (.sel({n172, n354, n181, n225}), .data({b[29], 
            1'b0, mulh[29], 1'bx}), .o(n859));   // alu.v(97)
    assign q1[29] = n849 ? n859 : 1'bz;   // alu.v(96)
    Select_4 Select_696 (.sel({n172, n354, n181, n225}), .data({b[28], 
            1'b0, mulh[28], 1'bx}), .o(n865));   // alu.v(97)
    assign q1[28] = n849 ? n865 : 1'bz;   // alu.v(96)
    Select_4 Select_702 (.sel({n172, n354, n181, n225}), .data({b[27], 
            1'b0, mulh[27], 1'bx}), .o(n871));   // alu.v(97)
    assign q1[27] = n849 ? n871 : 1'bz;   // alu.v(96)
    Select_4 Select_708 (.sel({n172, n354, n181, n225}), .data({b[26], 
            1'b0, mulh[26], 1'bx}), .o(n877));   // alu.v(97)
    assign q1[26] = n849 ? n877 : 1'bz;   // alu.v(96)
    Select_4 Select_714 (.sel({n172, n354, n181, n225}), .data({b[25], 
            1'b0, mulh[25], 1'bx}), .o(n883));   // alu.v(97)
    assign q1[25] = n849 ? n883 : 1'bz;   // alu.v(96)
    Select_4 Select_720 (.sel({n172, n354, n181, n225}), .data({b[24], 
            1'b0, mulh[24], 1'bx}), .o(n889));   // alu.v(97)
    assign q1[24] = n849 ? n889 : 1'bz;   // alu.v(96)
    Select_4 Select_726 (.sel({n172, n354, n181, n225}), .data({b[23], 
            1'b0, mulh[23], 1'bx}), .o(n895));   // alu.v(97)
    assign q1[23] = n849 ? n895 : 1'bz;   // alu.v(96)
    Select_4 Select_732 (.sel({n172, n354, n181, n225}), .data({b[22], 
            1'b0, mulh[22], 1'bx}), .o(n901));   // alu.v(97)
    assign q1[22] = n849 ? n901 : 1'bz;   // alu.v(96)
    Select_4 Select_738 (.sel({n172, n354, n181, n225}), .data({b[21], 
            1'b0, mulh[21], 1'bx}), .o(n907));   // alu.v(97)
    assign q1[21] = n849 ? n907 : 1'bz;   // alu.v(96)
    Select_4 Select_744 (.sel({n172, n354, n181, n225}), .data({b[20], 
            1'b0, mulh[20], 1'bx}), .o(n913));   // alu.v(97)
    assign q1[20] = n849 ? n913 : 1'bz;   // alu.v(96)
    Select_4 Select_750 (.sel({n172, n354, n181, n225}), .data({b[19], 
            1'b0, mulh[19], 1'bx}), .o(n919));   // alu.v(97)
    assign q1[19] = n849 ? n919 : 1'bz;   // alu.v(96)
    Select_4 Select_756 (.sel({n172, n354, n181, n225}), .data({b[18], 
            1'b0, mulh[18], 1'bx}), .o(n925));   // alu.v(97)
    assign q1[18] = n849 ? n925 : 1'bz;   // alu.v(96)
    Select_4 Select_762 (.sel({n172, n354, n181, n225}), .data({b[17], 
            1'b0, mulh[17], 1'bx}), .o(n931));   // alu.v(97)
    assign q1[17] = n849 ? n931 : 1'bz;   // alu.v(96)
    Select_4 Select_768 (.sel({n172, n354, n181, n225}), .data({b[16], 
            1'b0, mulh[16], 1'bx}), .o(n937));   // alu.v(97)
    assign q1[16] = n849 ? n937 : 1'bz;   // alu.v(96)
    Select_4 Select_774 (.sel({n172, n354, n181, n225}), .data({b[15], 
            1'b0, mulh[15], 1'bx}), .o(n943));   // alu.v(97)
    assign q1[15] = n849 ? n943 : 1'bz;   // alu.v(96)
    Select_4 Select_780 (.sel({n172, n354, n181, n225}), .data({b[14], 
            1'b0, mulh[14], 1'bx}), .o(n949));   // alu.v(97)
    assign q1[14] = n849 ? n949 : 1'bz;   // alu.v(96)
    Select_4 Select_786 (.sel({n172, n354, n181, n225}), .data({b[13], 
            1'b0, mulh[13], 1'bx}), .o(n955));   // alu.v(97)
    assign q1[13] = n849 ? n955 : 1'bz;   // alu.v(96)
    Select_4 Select_792 (.sel({n172, n354, n181, n225}), .data({b[12], 
            1'b0, mulh[12], 1'bx}), .o(n961));   // alu.v(97)
    assign q1[12] = n849 ? n961 : 1'bz;   // alu.v(96)
    Select_4 Select_798 (.sel({n172, n354, n181, n225}), .data({b[11], 
            1'b0, mulh[11], 1'bx}), .o(n967));   // alu.v(97)
    assign q1[11] = n849 ? n967 : 1'bz;   // alu.v(96)
    Select_4 Select_804 (.sel({n172, n354, n181, n225}), .data({b[10], 
            1'b0, mulh[10], 1'bx}), .o(n973));   // alu.v(97)
    assign q1[10] = n849 ? n973 : 1'bz;   // alu.v(96)
    Select_4 Select_810 (.sel({n172, n354, n181, n225}), .data({b[9], 
            1'b0, mulh[9], 1'bx}), .o(n979));   // alu.v(97)
    assign q1[9] = n849 ? n979 : 1'bz;   // alu.v(96)
    Select_4 Select_816 (.sel({n172, n354, n181, n225}), .data({b[8], 
            1'b0, mulh[8], 1'bx}), .o(n985));   // alu.v(97)
    assign q1[8] = n849 ? n985 : 1'bz;   // alu.v(96)
    Select_4 Select_822 (.sel({n172, n354, n181, n225}), .data({b[7], 
            1'b0, mulh[7], 1'bx}), .o(n991));   // alu.v(97)
    assign q1[7] = n849 ? n991 : 1'bz;   // alu.v(96)
    Select_4 Select_828 (.sel({n172, n354, n181, n225}), .data({b[6], 
            1'b0, mulh[6], 1'bx}), .o(n997));   // alu.v(97)
    assign q1[6] = n849 ? n997 : 1'bz;   // alu.v(96)
    Select_4 Select_834 (.sel({n172, n354, n181, n225}), .data({b[5], 
            1'b0, mulh[5], 1'bx}), .o(n1003));   // alu.v(97)
    assign q1[5] = n849 ? n1003 : 1'bz;   // alu.v(96)
    Select_4 Select_840 (.sel({n172, n354, n181, n225}), .data({b[4], 
            1'b0, mulh[4], 1'bx}), .o(n1009));   // alu.v(97)
    assign q1[4] = n849 ? n1009 : 1'bz;   // alu.v(96)
    Select_4 Select_846 (.sel({n172, n354, n181, n225}), .data({b[3], 
            1'b0, mulh[3], 1'bx}), .o(n1015));   // alu.v(97)
    assign q1[3] = n849 ? n1015 : 1'bz;   // alu.v(96)
    Select_4 Select_852 (.sel({n172, n354, n181, n225}), .data({b[2], 
            1'b0, mulh[2], 1'bx}), .o(n1021));   // alu.v(97)
    assign q1[2] = n849 ? n1021 : 1'bz;   // alu.v(96)
    Select_4 Select_858 (.sel({n172, n354, n181, n225}), .data({b[1], 
            1'b0, mulh[1], 1'bx}), .o(n1027));   // alu.v(97)
    assign q1[1] = n849 ? n1027 : 1'bz;   // alu.v(96)
    Select_4 Select_864 (.sel({n172, n354, n181, n225}), .data({b[0], 
            1'b0, mulh[0], 1'bx}), .o(n1033));   // alu.v(97)
    assign q1[0] = n849 ? n1033 : 1'bz;   // alu.v(96)
    Select_6 Select_870 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({1'b0, addsub[31], 1'b0, shift[31], 2'b0x}), .o(n1039));   // alu.v(97)
    assign st[3] = n657 ? n1039 : 1'bz;   // alu.v(96)
    Select_6 Select_876 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({1'b0, addsub_st[2], mul_st[2], shift_st[2], bws_st[2], 
            1'bx}), .o(n1045));   // alu.v(97)
    assign st[2] = n657 ? n1045 : 1'bz;   // alu.v(96)
    Select_6 Select_882 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({1'b0, addsub_st[1], mul_st[1], shift_st[1], 2'b0x}), 
            .o(n1051));   // alu.v(97)
    assign st[1] = n657 ? n1051 : 1'bz;   // alu.v(96)
    Select_6 Select_888 (.sel({n172, n226, n181, n227, n228, n225}), 
            .data({1'b0, addsub_st[0], 4'b000x}), .o(n1057));   // alu.v(97)
    assign st[0] = n657 ? n1057 : 1'bz;   // alu.v(96)
    Select_3 Select_894 (.sel({n434, n174, n435}), .data({3'bx01}), 
            .o(n1063));   // alu.v(97)
    Select_3 Select_896 (.sel({n434, n174, n435}), .data({3'b011}), 
            .o(n1065));   // alu.v(97)
    VERIFIC_DLATCHRS i904 (.d(n1069), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[31]));   // alu.v(96)
    Select_3 Select_900 (.sel({n434, n438, n179}), .data({1'bx, a[31], 
            1'b0}), .o(n1069));   // alu.v(97)
    Select_3 Select_902 (.sel({n434, n438, n179}), .data({3'b011}), 
            .o(n1071));   // alu.v(97)
    VERIFIC_DLATCHRS i910 (.d(n1075), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[30]));   // alu.v(96)
    Select_3 Select_906 (.sel({n434, n438, n179}), .data({1'bx, a[30], 
            1'b0}), .o(n1075));   // alu.v(97)
    VERIFIC_DLATCHRS i916 (.d(n1081), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[29]));   // alu.v(96)
    Select_3 Select_912 (.sel({n434, n438, n179}), .data({1'bx, a[29], 
            1'b0}), .o(n1081));   // alu.v(97)
    VERIFIC_DLATCHRS i922 (.d(n1087), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[28]));   // alu.v(96)
    Select_3 Select_918 (.sel({n434, n438, n179}), .data({1'bx, a[28], 
            1'b0}), .o(n1087));   // alu.v(97)
    VERIFIC_DLATCHRS i928 (.d(n1093), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[27]));   // alu.v(96)
    Select_3 Select_924 (.sel({n434, n438, n179}), .data({1'bx, a[27], 
            1'b0}), .o(n1093));   // alu.v(97)
    VERIFIC_DLATCHRS i934 (.d(n1099), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[26]));   // alu.v(96)
    Select_3 Select_930 (.sel({n434, n438, n179}), .data({1'bx, a[26], 
            1'b0}), .o(n1099));   // alu.v(97)
    VERIFIC_DLATCHRS i940 (.d(n1105), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[25]));   // alu.v(96)
    Select_3 Select_936 (.sel({n434, n438, n179}), .data({1'bx, a[25], 
            1'b0}), .o(n1105));   // alu.v(97)
    VERIFIC_DLATCHRS i946 (.d(n1111), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[24]));   // alu.v(96)
    Select_3 Select_942 (.sel({n434, n438, n179}), .data({1'bx, a[24], 
            1'b0}), .o(n1111));   // alu.v(97)
    VERIFIC_DLATCHRS i952 (.d(n1117), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[23]));   // alu.v(96)
    Select_3 Select_948 (.sel({n434, n438, n179}), .data({1'bx, a[23], 
            1'b0}), .o(n1117));   // alu.v(97)
    VERIFIC_DLATCHRS i958 (.d(n1123), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[22]));   // alu.v(96)
    Select_3 Select_954 (.sel({n434, n438, n179}), .data({1'bx, a[22], 
            1'b0}), .o(n1123));   // alu.v(97)
    VERIFIC_DLATCHRS i964 (.d(n1129), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[21]));   // alu.v(96)
    Select_3 Select_960 (.sel({n434, n438, n179}), .data({1'bx, a[21], 
            1'b0}), .o(n1129));   // alu.v(97)
    VERIFIC_DLATCHRS i970 (.d(n1135), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[20]));   // alu.v(96)
    Select_3 Select_966 (.sel({n434, n438, n179}), .data({1'bx, a[20], 
            1'b0}), .o(n1135));   // alu.v(97)
    VERIFIC_DLATCHRS i976 (.d(n1141), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[19]));   // alu.v(96)
    Select_3 Select_972 (.sel({n434, n438, n179}), .data({1'bx, a[19], 
            1'b0}), .o(n1141));   // alu.v(97)
    VERIFIC_DLATCHRS i982 (.d(n1147), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[18]));   // alu.v(96)
    Select_3 Select_978 (.sel({n434, n438, n179}), .data({1'bx, a[18], 
            1'b0}), .o(n1147));   // alu.v(97)
    VERIFIC_DLATCHRS i988 (.d(n1153), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[17]));   // alu.v(96)
    Select_3 Select_984 (.sel({n434, n438, n179}), .data({1'bx, a[17], 
            1'b0}), .o(n1153));   // alu.v(97)
    VERIFIC_DLATCHRS i994 (.d(n1159), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[16]));   // alu.v(96)
    Select_3 Select_990 (.sel({n434, n438, n179}), .data({1'bx, a[16], 
            1'b0}), .o(n1159));   // alu.v(97)
    VERIFIC_DLATCHRS i1000 (.d(n1165), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[15]));   // alu.v(96)
    Select_3 Select_996 (.sel({n434, n438, n179}), .data({1'bx, a[15], 
            1'b0}), .o(n1165));   // alu.v(97)
    VERIFIC_DLATCHRS i1006 (.d(n1171), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[14]));   // alu.v(96)
    Select_3 Select_1002 (.sel({n434, n438, n179}), .data({1'bx, a[14], 
            1'b0}), .o(n1171));   // alu.v(97)
    VERIFIC_DLATCHRS i1012 (.d(n1177), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[13]));   // alu.v(96)
    Select_3 Select_1008 (.sel({n434, n438, n179}), .data({1'bx, a[13], 
            1'b0}), .o(n1177));   // alu.v(97)
    VERIFIC_DLATCHRS i1018 (.d(n1183), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[12]));   // alu.v(96)
    Select_3 Select_1014 (.sel({n434, n438, n179}), .data({1'bx, a[12], 
            1'b0}), .o(n1183));   // alu.v(97)
    VERIFIC_DLATCHRS i1024 (.d(n1189), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[11]));   // alu.v(96)
    Select_3 Select_1020 (.sel({n434, n438, n179}), .data({1'bx, a[11], 
            1'b0}), .o(n1189));   // alu.v(97)
    VERIFIC_DLATCHRS i1030 (.d(n1195), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[10]));   // alu.v(96)
    Select_3 Select_1026 (.sel({n434, n438, n179}), .data({1'bx, a[10], 
            1'b0}), .o(n1195));   // alu.v(97)
    VERIFIC_DLATCHRS i1036 (.d(n1201), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[9]));   // alu.v(96)
    Select_3 Select_1032 (.sel({n434, n438, n179}), .data({1'bx, a[9], 
            1'b0}), .o(n1201));   // alu.v(97)
    VERIFIC_DLATCHRS i1042 (.d(n1207), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[8]));   // alu.v(96)
    Select_3 Select_1038 (.sel({n434, n438, n179}), .data({1'bx, a[8], 
            1'b0}), .o(n1207));   // alu.v(97)
    VERIFIC_DLATCHRS i1048 (.d(n1213), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[7]));   // alu.v(96)
    Select_3 Select_1044 (.sel({n434, n438, n179}), .data({1'bx, a[7], 
            1'b0}), .o(n1213));   // alu.v(97)
    VERIFIC_DLATCHRS i1054 (.d(n1219), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[6]));   // alu.v(96)
    Select_3 Select_1050 (.sel({n434, n438, n179}), .data({1'bx, a[6], 
            1'b0}), .o(n1219));   // alu.v(97)
    VERIFIC_DLATCHRS i1060 (.d(n1225), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[5]));   // alu.v(96)
    Select_3 Select_1056 (.sel({n434, n438, n179}), .data({1'bx, a[5], 
            1'b0}), .o(n1225));   // alu.v(97)
    VERIFIC_DLATCHRS i1066 (.d(n1231), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[4]));   // alu.v(96)
    Select_3 Select_1062 (.sel({n434, n438, n179}), .data({1'bx, a[4], 
            1'b0}), .o(n1231));   // alu.v(97)
    VERIFIC_DLATCHRS i1072 (.d(n1237), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[3]));   // alu.v(96)
    Select_3 Select_1068 (.sel({n434, n438, n179}), .data({1'bx, a[3], 
            1'b0}), .o(n1237));   // alu.v(97)
    VERIFIC_DLATCHRS i1078 (.d(n1243), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[2]));   // alu.v(96)
    Select_3 Select_1074 (.sel({n434, n438, n179}), .data({1'bx, a[2], 
            1'b0}), .o(n1243));   // alu.v(97)
    VERIFIC_DLATCHRS i1084 (.d(n1249), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[1]));   // alu.v(96)
    Select_3 Select_1080 (.sel({n434, n438, n179}), .data({1'bx, a[1], 
            1'b0}), .o(n1249));   // alu.v(97)
    VERIFIC_DLATCHRS i1090 (.d(n1255), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_a[0]));   // alu.v(96)
    Select_3 Select_1086 (.sel({n434, n438, n179}), .data({1'bx, a[0], 
            1'b0}), .o(n1255));   // alu.v(97)
    VERIFIC_DLATCHRS i1096 (.d(n1261), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[31]));   // alu.v(96)
    Select_3 Select_1092 (.sel({n434, n438, n179}), .data({1'bx, b[31], 
            a[31]}), .o(n1261));   // alu.v(97)
    VERIFIC_DLATCHRS i1102 (.d(n1267), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[30]));   // alu.v(96)
    Select_3 Select_1098 (.sel({n434, n438, n179}), .data({1'bx, b[30], 
            a[30]}), .o(n1267));   // alu.v(97)
    VERIFIC_DLATCHRS i1108 (.d(n1273), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[29]));   // alu.v(96)
    Select_3 Select_1104 (.sel({n434, n438, n179}), .data({1'bx, b[29], 
            a[29]}), .o(n1273));   // alu.v(97)
    VERIFIC_DLATCHRS i1114 (.d(n1279), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[28]));   // alu.v(96)
    Select_3 Select_1110 (.sel({n434, n438, n179}), .data({1'bx, b[28], 
            a[28]}), .o(n1279));   // alu.v(97)
    VERIFIC_DLATCHRS i1120 (.d(n1285), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[27]));   // alu.v(96)
    Select_3 Select_1116 (.sel({n434, n438, n179}), .data({1'bx, b[27], 
            a[27]}), .o(n1285));   // alu.v(97)
    VERIFIC_DLATCHRS i1126 (.d(n1291), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[26]));   // alu.v(96)
    Select_3 Select_1122 (.sel({n434, n438, n179}), .data({1'bx, b[26], 
            a[26]}), .o(n1291));   // alu.v(97)
    VERIFIC_DLATCHRS i1132 (.d(n1297), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[25]));   // alu.v(96)
    Select_3 Select_1128 (.sel({n434, n438, n179}), .data({1'bx, b[25], 
            a[25]}), .o(n1297));   // alu.v(97)
    VERIFIC_DLATCHRS i1138 (.d(n1303), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[24]));   // alu.v(96)
    Select_3 Select_1134 (.sel({n434, n438, n179}), .data({1'bx, b[24], 
            a[24]}), .o(n1303));   // alu.v(97)
    VERIFIC_DLATCHRS i1144 (.d(n1309), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[23]));   // alu.v(96)
    Select_3 Select_1140 (.sel({n434, n438, n179}), .data({1'bx, b[23], 
            a[23]}), .o(n1309));   // alu.v(97)
    VERIFIC_DLATCHRS i1150 (.d(n1315), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[22]));   // alu.v(96)
    Select_3 Select_1146 (.sel({n434, n438, n179}), .data({1'bx, b[22], 
            a[22]}), .o(n1315));   // alu.v(97)
    VERIFIC_DLATCHRS i1156 (.d(n1321), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[21]));   // alu.v(96)
    Select_3 Select_1152 (.sel({n434, n438, n179}), .data({1'bx, b[21], 
            a[21]}), .o(n1321));   // alu.v(97)
    VERIFIC_DLATCHRS i1162 (.d(n1327), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[20]));   // alu.v(96)
    Select_3 Select_1158 (.sel({n434, n438, n179}), .data({1'bx, b[20], 
            a[20]}), .o(n1327));   // alu.v(97)
    VERIFIC_DLATCHRS i1168 (.d(n1333), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[19]));   // alu.v(96)
    Select_3 Select_1164 (.sel({n434, n438, n179}), .data({1'bx, b[19], 
            a[19]}), .o(n1333));   // alu.v(97)
    VERIFIC_DLATCHRS i1174 (.d(n1339), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[18]));   // alu.v(96)
    Select_3 Select_1170 (.sel({n434, n438, n179}), .data({1'bx, b[18], 
            a[18]}), .o(n1339));   // alu.v(97)
    VERIFIC_DLATCHRS i1180 (.d(n1345), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[17]));   // alu.v(96)
    Select_3 Select_1176 (.sel({n434, n438, n179}), .data({1'bx, b[17], 
            a[17]}), .o(n1345));   // alu.v(97)
    VERIFIC_DLATCHRS i1186 (.d(n1351), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[16]));   // alu.v(96)
    Select_3 Select_1182 (.sel({n434, n438, n179}), .data({1'bx, b[16], 
            a[16]}), .o(n1351));   // alu.v(97)
    VERIFIC_DLATCHRS i1192 (.d(n1357), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[15]));   // alu.v(96)
    Select_3 Select_1188 (.sel({n434, n438, n179}), .data({1'bx, b[15], 
            a[15]}), .o(n1357));   // alu.v(97)
    VERIFIC_DLATCHRS i1198 (.d(n1363), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[14]));   // alu.v(96)
    Select_3 Select_1194 (.sel({n434, n438, n179}), .data({1'bx, b[14], 
            a[14]}), .o(n1363));   // alu.v(97)
    VERIFIC_DLATCHRS i1204 (.d(n1369), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[13]));   // alu.v(96)
    Select_3 Select_1200 (.sel({n434, n438, n179}), .data({1'bx, b[13], 
            a[13]}), .o(n1369));   // alu.v(97)
    VERIFIC_DLATCHRS i1210 (.d(n1375), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[12]));   // alu.v(96)
    Select_3 Select_1206 (.sel({n434, n438, n179}), .data({1'bx, b[12], 
            a[12]}), .o(n1375));   // alu.v(97)
    VERIFIC_DLATCHRS i1216 (.d(n1381), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[11]));   // alu.v(96)
    Select_3 Select_1212 (.sel({n434, n438, n179}), .data({1'bx, b[11], 
            a[11]}), .o(n1381));   // alu.v(97)
    VERIFIC_DLATCHRS i1222 (.d(n1387), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[10]));   // alu.v(96)
    Select_3 Select_1218 (.sel({n434, n438, n179}), .data({1'bx, b[10], 
            a[10]}), .o(n1387));   // alu.v(97)
    VERIFIC_DLATCHRS i1228 (.d(n1393), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[9]));   // alu.v(96)
    Select_3 Select_1224 (.sel({n434, n438, n179}), .data({1'bx, b[9], 
            a[9]}), .o(n1393));   // alu.v(97)
    VERIFIC_DLATCHRS i1234 (.d(n1399), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[8]));   // alu.v(96)
    Select_3 Select_1230 (.sel({n434, n438, n179}), .data({1'bx, b[8], 
            a[8]}), .o(n1399));   // alu.v(97)
    VERIFIC_DLATCHRS i1240 (.d(n1405), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[7]));   // alu.v(96)
    Select_3 Select_1236 (.sel({n434, n438, n179}), .data({1'bx, b[7], 
            a[7]}), .o(n1405));   // alu.v(97)
    VERIFIC_DLATCHRS i1246 (.d(n1411), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[6]));   // alu.v(96)
    Select_3 Select_1242 (.sel({n434, n438, n179}), .data({1'bx, b[6], 
            a[6]}), .o(n1411));   // alu.v(97)
    VERIFIC_DLATCHRS i1252 (.d(n1417), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[5]));   // alu.v(96)
    Select_3 Select_1248 (.sel({n434, n438, n179}), .data({1'bx, b[5], 
            a[5]}), .o(n1417));   // alu.v(97)
    VERIFIC_DLATCHRS i1258 (.d(n1423), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[4]));   // alu.v(96)
    Select_3 Select_1254 (.sel({n434, n438, n179}), .data({1'bx, b[4], 
            a[4]}), .o(n1423));   // alu.v(97)
    VERIFIC_DLATCHRS i1264 (.d(n1429), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[3]));   // alu.v(96)
    Select_3 Select_1260 (.sel({n434, n438, n179}), .data({1'bx, b[3], 
            a[3]}), .o(n1429));   // alu.v(97)
    VERIFIC_DLATCHRS i1270 (.d(n1435), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[2]));   // alu.v(96)
    Select_3 Select_1266 (.sel({n434, n438, n179}), .data({1'bx, b[2], 
            a[2]}), .o(n1435));   // alu.v(97)
    VERIFIC_DLATCHRS i1276 (.d(n1441), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[1]));   // alu.v(96)
    Select_3 Select_1272 (.sel({n434, n438, n179}), .data({1'bx, b[1], 
            a[1]}), .o(n1441));   // alu.v(97)
    VERIFIC_DLATCHRS i1282 (.d(n1447), .gate(n1071), .s(1'b0), .r(1'b0), 
            .q(addsub_b[0]));   // alu.v(96)
    Select_3 Select_1278 (.sel({n434, n438, n179}), .data({1'bx, b[0], 
            a[0]}), .o(n1447));   // alu.v(97)
    VERIFIC_DLATCHRS i1288 (.d(n1453), .gate(n1455), .s(1'b0), .r(1'b0), 
            .q(rotate));   // alu.v(96)
    Select_3 Select_1284 (.sel({n629, n630, n631}), .data({3'bx01}), 
            .o(n1453));   // alu.v(97)
    Select_3 Select_1286 (.sel({n629, n630, n631}), .data({3'b011}), 
            .o(n1455));   // alu.v(97)
    VERIFIC_DLATCHRS i1294 (.d(n1459), .gate(n1461), .s(1'b0), .r(1'b0), 
            .q(left));   // alu.v(96)
    Select_3 Select_1290 (.sel({n629, n634, n635}), .data({3'bx01}), 
            .o(n1459));   // alu.v(97)
    Select_3 Select_1292 (.sel({n629, n634, n635}), .data({3'b011}), 
            .o(n1461));   // alu.v(97)
    VERIFIC_DLATCHRS i1300 (.d(n1465), .gate(n1467), .s(1'b0), .r(1'b0), 
            .q(arithmetic));   // alu.v(96)
    Select_3 Select_1296 (.sel({n629, n638, n639}), .data({3'bx01}), 
            .o(n1465));   // alu.v(97)
    Select_3 Select_1298 (.sel({n629, n638, n639}), .data({3'b011}), 
            .o(n1467));   // alu.v(97)
    VERIFIC_DLATCHRS i1306 (.d(n1471), .gate(n1473), .s(1'b0), .r(1'b0), 
            .q(b_op[2]));   // alu.v(96)
    Select_3 Select_1302 (.sel({n641, n642, n643}), .data({3'bx01}), 
            .o(n1471));   // alu.v(97)
    Select_3 Select_1304 (.sel({n641, n642, n643}), .data({3'b011}), 
            .o(n1473));   // alu.v(97)
    VERIFIC_DLATCHRS i1312 (.d(n1477), .gate(n1479), .s(1'b0), .r(1'b0), 
            .q(b_op[1]));   // alu.v(96)
    Select_3 Select_1308 (.sel({n641, n646, n647}), .data({3'bx01}), 
            .o(n1477));   // alu.v(97)
    Select_3 Select_1310 (.sel({n641, n646, n647}), .data({3'b011}), 
            .o(n1479));   // alu.v(97)
    VERIFIC_DLATCHRS i1318 (.d(n1483), .gate(n1485), .s(1'b0), .r(1'b0), 
            .q(b_op[0]));   // alu.v(96)
    Select_3 Select_1314 (.sel({n641, n650, n651}), .data({3'bx01}), 
            .o(n1483));   // alu.v(97)
    Select_3 Select_1316 (.sel({n641, n650, n651}), .data({3'b011}), 
            .o(n1485));   // alu.v(97)
    VERIFIC_DLATCHRS i898 (.d(n1063), .gate(n1065), .s(1'b0), .r(1'b0), 
            .q(subtract));   // alu.v(96)
    
endmodule

//
// Verific Verilog Description of module addsub_32
//

module addsub_32 (q, a, b, sub, ov, sov, z);   // alu.v(6)
    output [31:0]q;   // alu.v(10)
    input [31:0]a;   // alu.v(7)
    input [31:0]b;   // alu.v(7)
    input sub;   // alu.v(8)
    output ov;   // alu.v(11)
    output sov;   // alu.v(11)
    output z;   // alu.v(11)
    
    wire [31:0]bm;   // alu.v(13)
    
    wire n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
        n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, 
        n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, 
        n35, n102, n104, n105, n106, n107;
    
    not (n4, b[31]) ;   // alu.v(13)
    not (n5, b[30]) ;   // alu.v(13)
    not (n6, b[29]) ;   // alu.v(13)
    not (n7, b[28]) ;   // alu.v(13)
    not (n8, b[27]) ;   // alu.v(13)
    not (n9, b[26]) ;   // alu.v(13)
    not (n10, b[25]) ;   // alu.v(13)
    not (n11, b[24]) ;   // alu.v(13)
    not (n12, b[23]) ;   // alu.v(13)
    not (n13, b[22]) ;   // alu.v(13)
    not (n14, b[21]) ;   // alu.v(13)
    not (n15, b[20]) ;   // alu.v(13)
    not (n16, b[19]) ;   // alu.v(13)
    not (n17, b[18]) ;   // alu.v(13)
    not (n18, b[17]) ;   // alu.v(13)
    not (n19, b[16]) ;   // alu.v(13)
    not (n20, b[15]) ;   // alu.v(13)
    not (n21, b[14]) ;   // alu.v(13)
    not (n22, b[13]) ;   // alu.v(13)
    not (n23, b[12]) ;   // alu.v(13)
    not (n24, b[11]) ;   // alu.v(13)
    not (n25, b[10]) ;   // alu.v(13)
    not (n26, b[9]) ;   // alu.v(13)
    not (n27, b[8]) ;   // alu.v(13)
    not (n28, b[7]) ;   // alu.v(13)
    not (n29, b[6]) ;   // alu.v(13)
    not (n30, b[5]) ;   // alu.v(13)
    not (n31, b[4]) ;   // alu.v(13)
    not (n32, b[3]) ;   // alu.v(13)
    not (n33, b[2]) ;   // alu.v(13)
    not (n34, b[1]) ;   // alu.v(13)
    not (n35, b[0]) ;   // alu.v(13)
    assign bm[31] = sub ? n4 : b[31];   // alu.v(13)
    assign bm[30] = sub ? n5 : b[30];   // alu.v(13)
    assign bm[29] = sub ? n6 : b[29];   // alu.v(13)
    assign bm[28] = sub ? n7 : b[28];   // alu.v(13)
    assign bm[27] = sub ? n8 : b[27];   // alu.v(13)
    assign bm[26] = sub ? n9 : b[26];   // alu.v(13)
    assign bm[25] = sub ? n10 : b[25];   // alu.v(13)
    assign bm[24] = sub ? n11 : b[24];   // alu.v(13)
    assign bm[23] = sub ? n12 : b[23];   // alu.v(13)
    assign bm[22] = sub ? n13 : b[22];   // alu.v(13)
    assign bm[21] = sub ? n14 : b[21];   // alu.v(13)
    assign bm[20] = sub ? n15 : b[20];   // alu.v(13)
    assign bm[19] = sub ? n16 : b[19];   // alu.v(13)
    assign bm[18] = sub ? n17 : b[18];   // alu.v(13)
    assign bm[17] = sub ? n18 : b[17];   // alu.v(13)
    assign bm[16] = sub ? n19 : b[16];   // alu.v(13)
    assign bm[15] = sub ? n20 : b[15];   // alu.v(13)
    assign bm[14] = sub ? n21 : b[14];   // alu.v(13)
    assign bm[13] = sub ? n22 : b[13];   // alu.v(13)
    assign bm[12] = sub ? n23 : b[12];   // alu.v(13)
    assign bm[11] = sub ? n24 : b[11];   // alu.v(13)
    assign bm[10] = sub ? n25 : b[10];   // alu.v(13)
    assign bm[9] = sub ? n26 : b[9];   // alu.v(13)
    assign bm[8] = sub ? n27 : b[8];   // alu.v(13)
    assign bm[7] = sub ? n28 : b[7];   // alu.v(13)
    assign bm[6] = sub ? n29 : b[6];   // alu.v(13)
    assign bm[5] = sub ? n30 : b[5];   // alu.v(13)
    assign bm[4] = sub ? n31 : b[4];   // alu.v(13)
    assign bm[3] = sub ? n32 : b[3];   // alu.v(13)
    assign bm[2] = sub ? n33 : b[2];   // alu.v(13)
    assign bm[1] = sub ? n34 : b[1];   // alu.v(13)
    assign bm[0] = sub ? n35 : b[0];   // alu.v(13)
    cla_32 cla0 (.a({a}), .b({bm}), .cin(sub), .s({q}), .cout(ov));   // alu.v(15)
    nor (z, q[31], q[30], q[29], q[28], q[27], q[26], q[25], 
           q[24], q[23], q[22], q[21], q[20], q[19], q[18], q[17], 
           q[16], q[15], q[14], q[13], q[12], q[11], q[10], q[9], 
           q[8], q[7], q[6], q[5], q[4], q[3], q[2], q[1], q[0]) ;   // alu.v(17)
    not (n102, a[31]) ;   // alu.v(19)
    and (n104, n102, n4) ;   // alu.v(19)
    and (n105, a[31], b[31]) ;   // alu.v(19)
    not (n106, q[31]) ;   // alu.v(19)
    assign n107 = n105 ? n106 : 1'b0;   // alu.v(19)
    assign sov = n104 ? ov : n107;   // alu.v(19)
    
endmodule

//
// Verific Verilog Description of module cla_32
//

module cla_32 (a, b, cin, s, cout);   // adder.v(70)
    input [31:0]a;   // adder.v(71)
    input [31:0]b;   // adder.v(72)
    input cin;   // adder.v(75)
    output [31:0]s;   // adder.v(73)
    output cout;   // adder.v(76)
    
    wire [3:0]p;   // adder.v(78)
    wire [3:0]g;   // adder.v(79)
    wire [2:0]c;   // adder.v(80)
    
    wire n40, n42, n43, n45;
    
    cla_16 cla0 (.a({a[15:0]}), .b({b[15:0]}), .cin(cin), .s({s[15:0]}), 
           .pg(p[0]), .gg(g[0]));   // adder.v(82)
    cla_16 cla1 (.a({a[31:16]}), .b({b[31:16]}), .cin(c[0]), .s({s[31:16]}), 
           .pg(p[1]), .gg(g[1]));   // adder.v(83)
    and (n40, p[0], cin) ;   // adder.v(85)
    or (c[0], g[0], n40) ;   // adder.v(85)
    and (n42, g[0], p[1]) ;   // adder.v(86)
    or (n43, g[1], n42) ;   // adder.v(86)
    and (n45, n40, p[1]) ;   // adder.v(86)
    or (cout, n43, n45) ;   // adder.v(86)
    
endmodule

//
// Verific Verilog Description of module cla_16
//

module cla_16 (a, b, cin, s, pg, gg);   // adder.v(44)
    input [15:0]a;   // adder.v(45)
    input [15:0]b;   // adder.v(46)
    input cin;   // adder.v(49)
    output [15:0]s;   // adder.v(47)
    output pg;   // adder.v(50)
    output gg;   // adder.v(50)
    
    wire [3:0]p;   // adder.v(52)
    wire [3:0]g;   // adder.v(53)
    wire [2:0]c;   // adder.v(54)
    
    wire n28, n30, n31, n33, n35, n36, n38, n39, n42, n44, 
        n45, n47, n48, n49, n50, n51, n52, n53, n54;
    
    cla_4 cla0 (.a({a[3:0]}), .b({b[3:0]}), .cin(cin), .s({s[3:0]}), 
          .pg(p[0]), .gg(g[0]));   // adder.v(56)
    cla_4 cla1 (.a({a[7:4]}), .b({b[7:4]}), .cin(c[0]), .s({s[7:4]}), 
          .pg(p[1]), .gg(g[1]));   // adder.v(57)
    cla_4 cla2 (.a({a[11:8]}), .b({b[11:8]}), .cin(c[1]), .s({s[11:8]}), 
          .pg(p[2]), .gg(g[2]));   // adder.v(58)
    cla_4 cla3 (.a({a[15:12]}), .b({b[15:12]}), .cin(c[2]), .s({s[15:12]}), 
          .pg(p[3]), .gg(g[3]));   // adder.v(59)
    and (n28, p[0], cin) ;   // adder.v(61)
    or (c[0], g[0], n28) ;   // adder.v(61)
    and (n30, g[0], p[1]) ;   // adder.v(62)
    or (n31, g[1], n30) ;   // adder.v(62)
    and (n33, n28, p[1]) ;   // adder.v(62)
    or (c[1], n31, n33) ;   // adder.v(62)
    and (n35, g[1], p[2]) ;   // adder.v(63)
    or (n36, g[2], n35) ;   // adder.v(63)
    and (n38, n30, p[2]) ;   // adder.v(63)
    or (n39, n36, n38) ;   // adder.v(63)
    and (n42, n33, p[2]) ;   // adder.v(63)
    or (c[2], n39, n42) ;   // adder.v(63)
    and (n44, p[0], p[1]) ;   // adder.v(65)
    and (n45, n44, p[2]) ;   // adder.v(65)
    and (pg, n45, p[3]) ;   // adder.v(65)
    and (n47, g[2], p[3]) ;   // adder.v(66)
    or (n48, g[3], n47) ;   // adder.v(66)
    and (n49, g[1], p[3]) ;   // adder.v(66)
    and (n50, n49, p[2]) ;   // adder.v(66)
    or (n51, n48, n50) ;   // adder.v(66)
    and (n52, g[0], p[3]) ;   // adder.v(66)
    and (n53, n52, p[2]) ;   // adder.v(66)
    and (n54, n53, p[1]) ;   // adder.v(66)
    or (gg, n51, n54) ;   // adder.v(66)
    
endmodule

//
// Verific Verilog Description of module cla_4
//

module cla_4 (a, b, cin, s, pg, gg);   // adder.v(18)
    input [3:0]a;   // adder.v(19)
    input [3:0]b;   // adder.v(20)
    input cin;   // adder.v(23)
    output [3:0]s;   // adder.v(21)
    output pg;   // adder.v(24)
    output gg;   // adder.v(24)
    
    wire [3:0]p;   // adder.v(26)
    wire [3:0]g;   // adder.v(27)
    wire [2:0]c;   // adder.v(28)
    
    wire n16, n18, n19, n21, n23, n24, n26, n27, n30, n32, 
        n33, n35, n36, n37, n38, n39, n40, n41, n42;
    
    fa_pg fa0 (.a(a[0]), .b(b[0]), .cin(cin), .s(s[0]), .p(p[0]), 
          .g(g[0]));   // adder.v(30)
    fa_pg fa1 (.a(a[1]), .b(b[1]), .cin(c[0]), .s(s[1]), .p(p[1]), 
          .g(g[1]));   // adder.v(31)
    fa_pg fa2 (.a(a[2]), .b(b[2]), .cin(c[1]), .s(s[2]), .p(p[2]), 
          .g(g[2]));   // adder.v(32)
    fa_pg fa3 (.a(a[3]), .b(b[3]), .cin(c[2]), .s(s[3]), .p(p[3]), 
          .g(g[3]));   // adder.v(33)
    and (n16, p[0], cin) ;   // adder.v(35)
    or (c[0], g[0], n16) ;   // adder.v(35)
    and (n18, g[0], p[1]) ;   // adder.v(36)
    or (n19, g[1], n18) ;   // adder.v(36)
    and (n21, n16, p[1]) ;   // adder.v(36)
    or (c[1], n19, n21) ;   // adder.v(36)
    and (n23, g[1], p[2]) ;   // adder.v(37)
    or (n24, g[2], n23) ;   // adder.v(37)
    and (n26, n18, p[2]) ;   // adder.v(37)
    or (n27, n24, n26) ;   // adder.v(37)
    and (n30, n21, p[2]) ;   // adder.v(37)
    or (c[2], n27, n30) ;   // adder.v(37)
    and (n32, p[0], p[1]) ;   // adder.v(39)
    and (n33, n32, p[2]) ;   // adder.v(39)
    and (pg, n33, p[3]) ;   // adder.v(39)
    and (n35, g[2], p[3]) ;   // adder.v(40)
    or (n36, g[3], n35) ;   // adder.v(40)
    and (n37, g[1], p[3]) ;   // adder.v(40)
    and (n38, n37, p[2]) ;   // adder.v(40)
    or (n39, n36, n38) ;   // adder.v(40)
    and (n40, g[0], p[3]) ;   // adder.v(40)
    and (n41, n40, p[2]) ;   // adder.v(40)
    and (n42, n41, p[1]) ;   // adder.v(40)
    or (gg, n39, n42) ;   // adder.v(40)
    
endmodule

//
// Verific Verilog Description of module fa_pg
//

module fa_pg (a, b, cin, s, p, g);   // adder.v(4)
    input a;   // adder.v(5)
    input b;   // adder.v(5)
    input cin;   // adder.v(5)
    output s;   // adder.v(7)
    output p;   // adder.v(7)
    output g;   // adder.v(7)
    
    
    xor (p, a, b) ;   // adder.v(11)
    xor (s, p, cin) ;   // adder.v(12)
    and (g, a, b) ;   // adder.v(14)
    
endmodule

//
// Verific Verilog Description of module bshift_32
//

module bshift_32 (q, ov, z, a, b, rotate, left, arith);   // shift.v(234)
    output [31:0]q;   // shift.v(239)
    output ov;   // shift.v(240)
    output z;   // shift.v(240)
    input [31:0]a;   // shift.v(235)
    input [4:0]b;   // shift.v(236)
    input rotate;   // shift.v(237)
    input left;   // shift.v(237)
    input arith;   // shift.v(237)
    
    wire [31:0]am;   // shift.v(242)
    wire [31:0]ym;   // shift.v(245)
    wire sra;   // shift.v(248)
    wire sla;   // shift.v(249)
    wire [31:0]f;   // shift.v(251)
    wire [31:0]p;   // shift.v(254)
    wire [31:0]t;   // shift.v(257)
    wire [31:0]zm;   // shift.v(262)
    
    wire n68, n69, n70, n73, n235, n236, n237, n238, n239, 
        n240, n241, n242, n243, n244, n245, n246, n247, n248, 
        n249, n250, n251, n252, n253, n254, n255, n256, n257, 
        n258, n259, n260, n261, n262, n263, n264, n265, n266;
    
    drev_32 dr0 (.q({am}), .a({a}), .e(left));   // shift.v(243)
    right_rot_32 rr0 (.y({ym}), .a({am}), .b({b}));   // shift.v(246)
    not (n68, rotate) ;   // shift.v(248)
    not (n69, left) ;   // shift.v(248)
    and (n70, n68, n69) ;   // shift.v(248)
    and (sra, n70, arith) ;   // shift.v(248)
    and (n73, n68, left) ;   // shift.v(249)
    and (sla, n73, arith) ;   // shift.v(249)
    fmask_32 f0 (.q({f}), .a({b}));   // shift.v(252)
    assign p[31] = rotate ? 1'b1 : f[31];   // shift.v(255)
    assign p[30] = rotate ? 1'b1 : f[30];   // shift.v(255)
    assign p[29] = rotate ? 1'b1 : f[29];   // shift.v(255)
    assign p[28] = rotate ? 1'b1 : f[28];   // shift.v(255)
    assign p[27] = rotate ? 1'b1 : f[27];   // shift.v(255)
    assign p[26] = rotate ? 1'b1 : f[26];   // shift.v(255)
    assign p[25] = rotate ? 1'b1 : f[25];   // shift.v(255)
    assign p[24] = rotate ? 1'b1 : f[24];   // shift.v(255)
    assign p[23] = rotate ? 1'b1 : f[23];   // shift.v(255)
    assign p[22] = rotate ? 1'b1 : f[22];   // shift.v(255)
    assign p[21] = rotate ? 1'b1 : f[21];   // shift.v(255)
    assign p[20] = rotate ? 1'b1 : f[20];   // shift.v(255)
    assign p[19] = rotate ? 1'b1 : f[19];   // shift.v(255)
    assign p[18] = rotate ? 1'b1 : f[18];   // shift.v(255)
    assign p[17] = rotate ? 1'b1 : f[17];   // shift.v(255)
    assign p[16] = rotate ? 1'b1 : f[16];   // shift.v(255)
    assign p[15] = rotate ? 1'b1 : f[15];   // shift.v(255)
    assign p[14] = rotate ? 1'b1 : f[14];   // shift.v(255)
    assign p[13] = rotate ? 1'b1 : f[13];   // shift.v(255)
    assign p[12] = rotate ? 1'b1 : f[12];   // shift.v(255)
    assign p[11] = rotate ? 1'b1 : f[11];   // shift.v(255)
    assign p[10] = rotate ? 1'b1 : f[10];   // shift.v(255)
    assign p[9] = rotate ? 1'b1 : f[9];   // shift.v(255)
    assign p[8] = rotate ? 1'b1 : f[8];   // shift.v(255)
    assign p[7] = rotate ? 1'b1 : f[7];   // shift.v(255)
    assign p[6] = rotate ? 1'b1 : f[6];   // shift.v(255)
    assign p[5] = rotate ? 1'b1 : f[5];   // shift.v(255)
    assign p[4] = rotate ? 1'b1 : f[4];   // shift.v(255)
    assign p[3] = rotate ? 1'b1 : f[3];   // shift.v(255)
    assign p[2] = rotate ? 1'b1 : f[2];   // shift.v(255)
    assign p[1] = rotate ? 1'b1 : f[1];   // shift.v(255)
    assign p[0] = rotate ? 1'b1 : f[0];   // shift.v(255)
    tblock_32 t0 (.q({t}), .a({ym}), .sgn(a[31]), .p({p}), .sla(sla), 
            .sra(sra));   // shift.v(258)
    drev_32 dr1 (.q({q}), .a({t}), .e(left));   // shift.v(260)
    zmask_32 z0 (.q({zm}), .a({p}), .sla(sla));   // shift.v(263)
    and (n235, zm[0], am[0]) ;   // shift.v(265)
    and (n236, zm[1], am[1]) ;   // shift.v(265)
    and (n237, zm[2], am[2]) ;   // shift.v(265)
    and (n238, zm[3], am[3]) ;   // shift.v(265)
    and (n239, zm[4], am[4]) ;   // shift.v(265)
    and (n240, zm[5], am[5]) ;   // shift.v(265)
    and (n241, zm[6], am[6]) ;   // shift.v(265)
    and (n242, zm[7], am[7]) ;   // shift.v(265)
    and (n243, zm[8], am[8]) ;   // shift.v(265)
    and (n244, zm[9], am[9]) ;   // shift.v(265)
    and (n245, zm[10], am[10]) ;   // shift.v(265)
    and (n246, zm[11], am[11]) ;   // shift.v(265)
    and (n247, zm[12], am[12]) ;   // shift.v(265)
    and (n248, zm[13], am[13]) ;   // shift.v(265)
    and (n249, zm[14], am[14]) ;   // shift.v(265)
    and (n250, zm[15], am[15]) ;   // shift.v(265)
    and (n251, zm[16], am[16]) ;   // shift.v(265)
    and (n252, zm[17], am[17]) ;   // shift.v(265)
    and (n253, zm[18], am[18]) ;   // shift.v(265)
    and (n254, zm[19], am[19]) ;   // shift.v(265)
    and (n255, zm[20], am[20]) ;   // shift.v(265)
    and (n256, zm[21], am[21]) ;   // shift.v(265)
    and (n257, zm[22], am[22]) ;   // shift.v(265)
    and (n258, zm[23], am[23]) ;   // shift.v(265)
    and (n259, zm[24], am[24]) ;   // shift.v(265)
    and (n260, zm[25], am[25]) ;   // shift.v(265)
    and (n261, zm[26], am[26]) ;   // shift.v(265)
    and (n262, zm[27], am[27]) ;   // shift.v(265)
    and (n263, zm[28], am[28]) ;   // shift.v(265)
    and (n264, zm[29], am[29]) ;   // shift.v(265)
    and (n265, zm[30], am[30]) ;   // shift.v(265)
    and (n266, zm[31], am[31]) ;   // shift.v(265)
    nor (z, n266, n265, n264, n263, n262, n261, n260, n259, 
        n258, n257, n256, n255, n254, n253, n252, n251, n250, 
        n249, n248, n247, n246, n245, n244, n243, n242, n241, 
        n240, n239, n238, n237, n236, n235) ;   // shift.v(265)
    ovf_32 ov0 (.q(ov), .a({a}), .f({f}), .sla(sla));   // shift.v(267)
    
endmodule

//
// Verific Verilog Description of module drev_32
//

module drev_32 (q, a, e);   // shift.v(135)
    output [31:0]q;   // shift.v(138)
    input [31:0]a;   // shift.v(136)
    input e;   // shift.v(139)
    
    
    assign q[0] = e ? a[31] : a[0];   // shift.v(143)
    assign q[1] = e ? a[30] : a[1];   // shift.v(143)
    assign q[2] = e ? a[29] : a[2];   // shift.v(143)
    assign q[3] = e ? a[28] : a[3];   // shift.v(143)
    assign q[4] = e ? a[27] : a[4];   // shift.v(143)
    assign q[5] = e ? a[26] : a[5];   // shift.v(143)
    assign q[6] = e ? a[25] : a[6];   // shift.v(143)
    assign q[7] = e ? a[24] : a[7];   // shift.v(143)
    assign q[8] = e ? a[23] : a[8];   // shift.v(143)
    assign q[9] = e ? a[22] : a[9];   // shift.v(143)
    assign q[10] = e ? a[21] : a[10];   // shift.v(143)
    assign q[11] = e ? a[20] : a[11];   // shift.v(143)
    assign q[12] = e ? a[19] : a[12];   // shift.v(143)
    assign q[13] = e ? a[18] : a[13];   // shift.v(143)
    assign q[14] = e ? a[17] : a[14];   // shift.v(143)
    assign q[15] = e ? a[16] : a[15];   // shift.v(143)
    assign q[16] = e ? a[15] : a[16];   // shift.v(143)
    assign q[17] = e ? a[14] : a[17];   // shift.v(143)
    assign q[18] = e ? a[13] : a[18];   // shift.v(143)
    assign q[19] = e ? a[12] : a[19];   // shift.v(143)
    assign q[20] = e ? a[11] : a[20];   // shift.v(143)
    assign q[21] = e ? a[10] : a[21];   // shift.v(143)
    assign q[22] = e ? a[9] : a[22];   // shift.v(143)
    assign q[23] = e ? a[8] : a[23];   // shift.v(143)
    assign q[24] = e ? a[7] : a[24];   // shift.v(143)
    assign q[25] = e ? a[6] : a[25];   // shift.v(143)
    assign q[26] = e ? a[5] : a[26];   // shift.v(143)
    assign q[27] = e ? a[4] : a[27];   // shift.v(143)
    assign q[28] = e ? a[3] : a[28];   // shift.v(143)
    assign q[29] = e ? a[2] : a[29];   // shift.v(143)
    assign q[30] = e ? a[1] : a[30];   // shift.v(143)
    assign q[31] = e ? a[0] : a[31];   // shift.v(143)
    
endmodule

//
// Verific Verilog Description of module right_rot_32
//

module right_rot_32 (y, a, b);   // shift.v(103)
    output [31:0]y;   // shift.v(107)
    input [31:0]a;   // shift.v(104)
    input [4:0]b;   // shift.v(105)
    
    wire [31:0]st1;   // shift.v(110)
    wire [31:0]st2;   // shift.v(115)
    wire [31:0]st3;   // shift.v(120)
    wire [31:0]st4;   // shift.v(125)
    
    assign st1[31] = b[4] ? a[15] : a[31];   // shift.v(112)
    assign st1[30] = b[4] ? a[14] : a[30];   // shift.v(112)
    assign st1[29] = b[4] ? a[13] : a[29];   // shift.v(112)
    assign st1[28] = b[4] ? a[12] : a[28];   // shift.v(112)
    assign st1[27] = b[4] ? a[11] : a[27];   // shift.v(112)
    assign st1[26] = b[4] ? a[10] : a[26];   // shift.v(112)
    assign st1[25] = b[4] ? a[9] : a[25];   // shift.v(112)
    assign st1[24] = b[4] ? a[8] : a[24];   // shift.v(112)
    assign st1[23] = b[4] ? a[7] : a[23];   // shift.v(112)
    assign st1[22] = b[4] ? a[6] : a[22];   // shift.v(112)
    assign st1[21] = b[4] ? a[5] : a[21];   // shift.v(112)
    assign st1[20] = b[4] ? a[4] : a[20];   // shift.v(112)
    assign st1[19] = b[4] ? a[3] : a[19];   // shift.v(112)
    assign st1[18] = b[4] ? a[2] : a[18];   // shift.v(112)
    assign st1[17] = b[4] ? a[1] : a[17];   // shift.v(112)
    assign st1[16] = b[4] ? a[0] : a[16];   // shift.v(112)
    assign st1[15] = b[4] ? a[31] : a[15];   // shift.v(113)
    assign st1[14] = b[4] ? a[30] : a[14];   // shift.v(113)
    assign st1[13] = b[4] ? a[29] : a[13];   // shift.v(113)
    assign st1[12] = b[4] ? a[28] : a[12];   // shift.v(113)
    assign st1[11] = b[4] ? a[27] : a[11];   // shift.v(113)
    assign st1[10] = b[4] ? a[26] : a[10];   // shift.v(113)
    assign st1[9] = b[4] ? a[25] : a[9];   // shift.v(113)
    assign st1[8] = b[4] ? a[24] : a[8];   // shift.v(113)
    assign st1[7] = b[4] ? a[23] : a[7];   // shift.v(113)
    assign st1[6] = b[4] ? a[22] : a[6];   // shift.v(113)
    assign st1[5] = b[4] ? a[21] : a[5];   // shift.v(113)
    assign st1[4] = b[4] ? a[20] : a[4];   // shift.v(113)
    assign st1[3] = b[4] ? a[19] : a[3];   // shift.v(113)
    assign st1[2] = b[4] ? a[18] : a[2];   // shift.v(113)
    assign st1[1] = b[4] ? a[17] : a[1];   // shift.v(113)
    assign st1[0] = b[4] ? a[16] : a[0];   // shift.v(113)
    assign st2[31] = b[3] ? st1[7] : st1[31];   // shift.v(117)
    assign st2[30] = b[3] ? st1[6] : st1[30];   // shift.v(117)
    assign st2[29] = b[3] ? st1[5] : st1[29];   // shift.v(117)
    assign st2[28] = b[3] ? st1[4] : st1[28];   // shift.v(117)
    assign st2[27] = b[3] ? st1[3] : st1[27];   // shift.v(117)
    assign st2[26] = b[3] ? st1[2] : st1[26];   // shift.v(117)
    assign st2[25] = b[3] ? st1[1] : st1[25];   // shift.v(117)
    assign st2[24] = b[3] ? st1[0] : st1[24];   // shift.v(117)
    assign st2[23] = b[3] ? st1[31] : st1[23];   // shift.v(118)
    assign st2[22] = b[3] ? st1[30] : st1[22];   // shift.v(118)
    assign st2[21] = b[3] ? st1[29] : st1[21];   // shift.v(118)
    assign st2[20] = b[3] ? st1[28] : st1[20];   // shift.v(118)
    assign st2[19] = b[3] ? st1[27] : st1[19];   // shift.v(118)
    assign st2[18] = b[3] ? st1[26] : st1[18];   // shift.v(118)
    assign st2[17] = b[3] ? st1[25] : st1[17];   // shift.v(118)
    assign st2[16] = b[3] ? st1[24] : st1[16];   // shift.v(118)
    assign st2[15] = b[3] ? st1[23] : st1[15];   // shift.v(118)
    assign st2[14] = b[3] ? st1[22] : st1[14];   // shift.v(118)
    assign st2[13] = b[3] ? st1[21] : st1[13];   // shift.v(118)
    assign st2[12] = b[3] ? st1[20] : st1[12];   // shift.v(118)
    assign st2[11] = b[3] ? st1[19] : st1[11];   // shift.v(118)
    assign st2[10] = b[3] ? st1[18] : st1[10];   // shift.v(118)
    assign st2[9] = b[3] ? st1[17] : st1[9];   // shift.v(118)
    assign st2[8] = b[3] ? st1[16] : st1[8];   // shift.v(118)
    assign st2[7] = b[3] ? st1[15] : st1[7];   // shift.v(118)
    assign st2[6] = b[3] ? st1[14] : st1[6];   // shift.v(118)
    assign st2[5] = b[3] ? st1[13] : st1[5];   // shift.v(118)
    assign st2[4] = b[3] ? st1[12] : st1[4];   // shift.v(118)
    assign st2[3] = b[3] ? st1[11] : st1[3];   // shift.v(118)
    assign st2[2] = b[3] ? st1[10] : st1[2];   // shift.v(118)
    assign st2[1] = b[3] ? st1[9] : st1[1];   // shift.v(118)
    assign st2[0] = b[3] ? st1[8] : st1[0];   // shift.v(118)
    assign st3[31] = b[2] ? st2[3] : st2[31];   // shift.v(122)
    assign st3[30] = b[2] ? st2[2] : st2[30];   // shift.v(122)
    assign st3[29] = b[2] ? st2[1] : st2[29];   // shift.v(122)
    assign st3[28] = b[2] ? st2[0] : st2[28];   // shift.v(122)
    assign st3[27] = b[2] ? st2[31] : st2[27];   // shift.v(123)
    assign st3[26] = b[2] ? st2[30] : st2[26];   // shift.v(123)
    assign st3[25] = b[2] ? st2[29] : st2[25];   // shift.v(123)
    assign st3[24] = b[2] ? st2[28] : st2[24];   // shift.v(123)
    assign st3[23] = b[2] ? st2[27] : st2[23];   // shift.v(123)
    assign st3[22] = b[2] ? st2[26] : st2[22];   // shift.v(123)
    assign st3[21] = b[2] ? st2[25] : st2[21];   // shift.v(123)
    assign st3[20] = b[2] ? st2[24] : st2[20];   // shift.v(123)
    assign st3[19] = b[2] ? st2[23] : st2[19];   // shift.v(123)
    assign st3[18] = b[2] ? st2[22] : st2[18];   // shift.v(123)
    assign st3[17] = b[2] ? st2[21] : st2[17];   // shift.v(123)
    assign st3[16] = b[2] ? st2[20] : st2[16];   // shift.v(123)
    assign st3[15] = b[2] ? st2[19] : st2[15];   // shift.v(123)
    assign st3[14] = b[2] ? st2[18] : st2[14];   // shift.v(123)
    assign st3[13] = b[2] ? st2[17] : st2[13];   // shift.v(123)
    assign st3[12] = b[2] ? st2[16] : st2[12];   // shift.v(123)
    assign st3[11] = b[2] ? st2[15] : st2[11];   // shift.v(123)
    assign st3[10] = b[2] ? st2[14] : st2[10];   // shift.v(123)
    assign st3[9] = b[2] ? st2[13] : st2[9];   // shift.v(123)
    assign st3[8] = b[2] ? st2[12] : st2[8];   // shift.v(123)
    assign st3[7] = b[2] ? st2[11] : st2[7];   // shift.v(123)
    assign st3[6] = b[2] ? st2[10] : st2[6];   // shift.v(123)
    assign st3[5] = b[2] ? st2[9] : st2[5];   // shift.v(123)
    assign st3[4] = b[2] ? st2[8] : st2[4];   // shift.v(123)
    assign st3[3] = b[2] ? st2[7] : st2[3];   // shift.v(123)
    assign st3[2] = b[2] ? st2[6] : st2[2];   // shift.v(123)
    assign st3[1] = b[2] ? st2[5] : st2[1];   // shift.v(123)
    assign st3[0] = b[2] ? st2[4] : st2[0];   // shift.v(123)
    assign st4[31] = b[1] ? st3[1] : st3[31];   // shift.v(127)
    assign st4[30] = b[1] ? st3[0] : st3[30];   // shift.v(127)
    assign st4[29] = b[1] ? st3[31] : st3[29];   // shift.v(128)
    assign st4[28] = b[1] ? st3[30] : st3[28];   // shift.v(128)
    assign st4[27] = b[1] ? st3[29] : st3[27];   // shift.v(128)
    assign st4[26] = b[1] ? st3[28] : st3[26];   // shift.v(128)
    assign st4[25] = b[1] ? st3[27] : st3[25];   // shift.v(128)
    assign st4[24] = b[1] ? st3[26] : st3[24];   // shift.v(128)
    assign st4[23] = b[1] ? st3[25] : st3[23];   // shift.v(128)
    assign st4[22] = b[1] ? st3[24] : st3[22];   // shift.v(128)
    assign st4[21] = b[1] ? st3[23] : st3[21];   // shift.v(128)
    assign st4[20] = b[1] ? st3[22] : st3[20];   // shift.v(128)
    assign st4[19] = b[1] ? st3[21] : st3[19];   // shift.v(128)
    assign st4[18] = b[1] ? st3[20] : st3[18];   // shift.v(128)
    assign st4[17] = b[1] ? st3[19] : st3[17];   // shift.v(128)
    assign st4[16] = b[1] ? st3[18] : st3[16];   // shift.v(128)
    assign st4[15] = b[1] ? st3[17] : st3[15];   // shift.v(128)
    assign st4[14] = b[1] ? st3[16] : st3[14];   // shift.v(128)
    assign st4[13] = b[1] ? st3[15] : st3[13];   // shift.v(128)
    assign st4[12] = b[1] ? st3[14] : st3[12];   // shift.v(128)
    assign st4[11] = b[1] ? st3[13] : st3[11];   // shift.v(128)
    assign st4[10] = b[1] ? st3[12] : st3[10];   // shift.v(128)
    assign st4[9] = b[1] ? st3[11] : st3[9];   // shift.v(128)
    assign st4[8] = b[1] ? st3[10] : st3[8];   // shift.v(128)
    assign st4[7] = b[1] ? st3[9] : st3[7];   // shift.v(128)
    assign st4[6] = b[1] ? st3[8] : st3[6];   // shift.v(128)
    assign st4[5] = b[1] ? st3[7] : st3[5];   // shift.v(128)
    assign st4[4] = b[1] ? st3[6] : st3[4];   // shift.v(128)
    assign st4[3] = b[1] ? st3[5] : st3[3];   // shift.v(128)
    assign st4[2] = b[1] ? st3[4] : st3[2];   // shift.v(128)
    assign st4[1] = b[1] ? st3[3] : st3[1];   // shift.v(128)
    assign st4[0] = b[1] ? st3[2] : st3[0];   // shift.v(128)
    assign y[31] = b[0] ? st4[0] : st4[31];   // shift.v(131)
    assign y[30] = b[0] ? st4[31] : st4[30];   // shift.v(132)
    assign y[29] = b[0] ? st4[30] : st4[29];   // shift.v(132)
    assign y[28] = b[0] ? st4[29] : st4[28];   // shift.v(132)
    assign y[27] = b[0] ? st4[28] : st4[27];   // shift.v(132)
    assign y[26] = b[0] ? st4[27] : st4[26];   // shift.v(132)
    assign y[25] = b[0] ? st4[26] : st4[25];   // shift.v(132)
    assign y[24] = b[0] ? st4[25] : st4[24];   // shift.v(132)
    assign y[23] = b[0] ? st4[24] : st4[23];   // shift.v(132)
    assign y[22] = b[0] ? st4[23] : st4[22];   // shift.v(132)
    assign y[21] = b[0] ? st4[22] : st4[21];   // shift.v(132)
    assign y[20] = b[0] ? st4[21] : st4[20];   // shift.v(132)
    assign y[19] = b[0] ? st4[20] : st4[19];   // shift.v(132)
    assign y[18] = b[0] ? st4[19] : st4[18];   // shift.v(132)
    assign y[17] = b[0] ? st4[18] : st4[17];   // shift.v(132)
    assign y[16] = b[0] ? st4[17] : st4[16];   // shift.v(132)
    assign y[15] = b[0] ? st4[16] : st4[15];   // shift.v(132)
    assign y[14] = b[0] ? st4[15] : st4[14];   // shift.v(132)
    assign y[13] = b[0] ? st4[14] : st4[13];   // shift.v(132)
    assign y[12] = b[0] ? st4[13] : st4[12];   // shift.v(132)
    assign y[11] = b[0] ? st4[12] : st4[11];   // shift.v(132)
    assign y[10] = b[0] ? st4[11] : st4[10];   // shift.v(132)
    assign y[9] = b[0] ? st4[10] : st4[9];   // shift.v(132)
    assign y[8] = b[0] ? st4[9] : st4[8];   // shift.v(132)
    assign y[7] = b[0] ? st4[8] : st4[7];   // shift.v(132)
    assign y[6] = b[0] ? st4[7] : st4[6];   // shift.v(132)
    assign y[5] = b[0] ? st4[6] : st4[5];   // shift.v(132)
    assign y[4] = b[0] ? st4[5] : st4[4];   // shift.v(132)
    assign y[3] = b[0] ? st4[4] : st4[3];   // shift.v(132)
    assign y[2] = b[0] ? st4[3] : st4[2];   // shift.v(132)
    assign y[1] = b[0] ? st4[2] : st4[1];   // shift.v(132)
    assign y[0] = b[0] ? st4[1] : st4[0];   // shift.v(132)
    
endmodule

//
// Verific Verilog Description of module fmask_32
//

module fmask_32 (q, a);   // shift.v(148)
    output [31:0]q;   // shift.v(150)
    input [4:0]a;   // shift.v(149)
    
    
    assign q[0] = 1'b1;
    Mux_5u_32u Mux_3 (.sel({a}), .data({32'b00000000000000000000000000000001}), 
            .o(q[31]));   // shift.v(154)
    Mux_4u_16u Mux_4 (.sel({a[4:1]}), .data({16'b0000000000000001}), .o(q[30]));   // shift.v(154)
    Mux_5u_32u Mux_5 (.sel({a}), .data({32'b00000000000000000000000000000111}), 
            .o(q[29]));   // shift.v(154)
    Mux_3u_8u Mux_6 (.sel({a[4:2]}), .data({8'b00000001}), .o(q[28]));   // shift.v(154)
    Mux_5u_32u Mux_7 (.sel({a}), .data({32'b00000000000000000000000000011111}), 
            .o(q[27]));   // shift.v(154)
    Mux_4u_16u Mux_8 (.sel({a[4:1]}), .data({16'b0000000000000111}), .o(q[26]));   // shift.v(154)
    Mux_5u_32u Mux_9 (.sel({a}), .data({32'b00000000000000000000000001111111}), 
            .o(q[25]));   // shift.v(154)
    Mux_2u_4u Mux_10 (.sel({a[4:3]}), .data({4'b0001}), .o(q[24]));   // shift.v(154)
    Mux_5u_32u Mux_11 (.sel({a}), .data({32'b00000000000000000000000111111111}), 
            .o(q[23]));   // shift.v(154)
    Mux_4u_16u Mux_12 (.sel({a[4:1]}), .data({16'b0000000000011111}), .o(q[22]));   // shift.v(154)
    Mux_5u_32u Mux_13 (.sel({a}), .data({32'b00000000000000000000011111111111}), 
            .o(q[21]));   // shift.v(154)
    Mux_3u_8u Mux_14 (.sel({a[4:2]}), .data({8'b00000111}), .o(q[20]));   // shift.v(154)
    Mux_5u_32u Mux_15 (.sel({a}), .data({32'b00000000000000000001111111111111}), 
            .o(q[19]));   // shift.v(154)
    Mux_4u_16u Mux_16 (.sel({a[4:1]}), .data({16'b0000000001111111}), .o(q[18]));   // shift.v(154)
    Mux_5u_32u Mux_17 (.sel({a}), .data({32'b00000000000000000111111111111111}), 
            .o(q[17]));   // shift.v(154)
    not (q[16], a[4]) ;   // shift.v(154)
    Mux_5u_32u Mux_19 (.sel({a}), .data({32'b00000000000000011111111111111111}), 
            .o(q[15]));   // shift.v(154)
    Mux_4u_16u Mux_20 (.sel({a[4:1]}), .data({16'b0000000111111111}), .o(q[14]));   // shift.v(154)
    Mux_5u_32u Mux_21 (.sel({a}), .data({32'b00000000000001111111111111111111}), 
            .o(q[13]));   // shift.v(154)
    Mux_3u_8u Mux_22 (.sel({a[4:2]}), .data({8'b00011111}), .o(q[12]));   // shift.v(154)
    Mux_5u_32u Mux_23 (.sel({a}), .data({32'b00000000000111111111111111111111}), 
            .o(q[11]));   // shift.v(154)
    Mux_4u_16u Mux_24 (.sel({a[4:1]}), .data({16'b0000011111111111}), .o(q[10]));   // shift.v(154)
    Mux_5u_32u Mux_25 (.sel({a}), .data({32'b00000000011111111111111111111111}), 
            .o(q[9]));   // shift.v(154)
    Mux_2u_4u Mux_26 (.sel({a[4:3]}), .data({4'b0111}), .o(q[8]));   // shift.v(154)
    Mux_5u_32u Mux_27 (.sel({a}), .data({32'b00000001111111111111111111111111}), 
            .o(q[7]));   // shift.v(154)
    Mux_4u_16u Mux_28 (.sel({a[4:1]}), .data({16'b0001111111111111}), .o(q[6]));   // shift.v(154)
    Mux_5u_32u Mux_29 (.sel({a}), .data({32'b00000111111111111111111111111111}), 
            .o(q[5]));   // shift.v(154)
    Mux_3u_8u Mux_30 (.sel({a[4:2]}), .data({8'b01111111}), .o(q[4]));   // shift.v(154)
    Mux_5u_32u Mux_31 (.sel({a}), .data({32'b00011111111111111111111111111111}), 
            .o(q[3]));   // shift.v(154)
    Mux_4u_16u Mux_32 (.sel({a[4:1]}), .data({16'b0111111111111111}), .o(q[2]));   // shift.v(154)
    Mux_5u_32u Mux_33 (.sel({a}), .data({32'b01111111111111111111111111111111}), 
            .o(q[1]));   // shift.v(154)
    
endmodule

//
// Verific Verilog Description of OPERATOR Mux_4u_16u
//

module Mux_4u_16u (sel, data, o);
    input [3:0]sel;
    input [15:0]data;
    output o;
    assign o = data[sel];
    
endmodule

//
// Verific Verilog Description of OPERATOR Mux_3u_8u
//

module Mux_3u_8u (sel, data, o);
    input [2:0]sel;
    input [7:0]data;
    output o;
    assign o = data[sel];
    
endmodule

//
// Verific Verilog Description of OPERATOR Mux_2u_4u
//

module Mux_2u_4u (sel, data, o);
    input [1:0]sel;
    input [3:0]data;
    output o;
    assign o = data[sel];
    
endmodule

//
// Verific Verilog Description of module tblock_32
//

module tblock_32 (q, a, sgn, p, sla, sra);   // shift.v(221)
    output [31:0]q;   // shift.v(226)
    input [31:0]a;   // shift.v(222)
    input sgn;   // shift.v(224)
    input [31:0]p;   // shift.v(223)
    input sla;   // shift.v(224)
    input sra;   // shift.v(224)
    
    wire [30:0]s;   // shift.v(228)
    
    wire n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, 
        n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, 
        n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, 
        n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
        n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, 
        n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
        n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
        n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, 
        n97, n98, n99, n100, n101;
    
    and (s[30], sra, sgn) ;   // shift.v(228)
    not (n5, sla) ;   // shift.v(230)
    and (n6, a[0], n5) ;   // shift.v(230)
    and (n7, sla, sgn) ;   // shift.v(230)
    or (q[0], n6, n7) ;   // shift.v(230)
    and (n9, a[1], p[1]) ;   // shift.v(231)
    and (n10, a[2], p[2]) ;   // shift.v(231)
    and (n11, a[3], p[3]) ;   // shift.v(231)
    and (n12, a[4], p[4]) ;   // shift.v(231)
    and (n13, a[5], p[5]) ;   // shift.v(231)
    and (n14, a[6], p[6]) ;   // shift.v(231)
    and (n15, a[7], p[7]) ;   // shift.v(231)
    and (n16, a[8], p[8]) ;   // shift.v(231)
    and (n17, a[9], p[9]) ;   // shift.v(231)
    and (n18, a[10], p[10]) ;   // shift.v(231)
    and (n19, a[11], p[11]) ;   // shift.v(231)
    and (n20, a[12], p[12]) ;   // shift.v(231)
    and (n21, a[13], p[13]) ;   // shift.v(231)
    and (n22, a[14], p[14]) ;   // shift.v(231)
    and (n23, a[15], p[15]) ;   // shift.v(231)
    and (n24, a[16], p[16]) ;   // shift.v(231)
    and (n25, a[17], p[17]) ;   // shift.v(231)
    and (n26, a[18], p[18]) ;   // shift.v(231)
    and (n27, a[19], p[19]) ;   // shift.v(231)
    and (n28, a[20], p[20]) ;   // shift.v(231)
    and (n29, a[21], p[21]) ;   // shift.v(231)
    and (n30, a[22], p[22]) ;   // shift.v(231)
    and (n31, a[23], p[23]) ;   // shift.v(231)
    and (n32, a[24], p[24]) ;   // shift.v(231)
    and (n33, a[25], p[25]) ;   // shift.v(231)
    and (n34, a[26], p[26]) ;   // shift.v(231)
    and (n35, a[27], p[27]) ;   // shift.v(231)
    and (n36, a[28], p[28]) ;   // shift.v(231)
    and (n37, a[29], p[29]) ;   // shift.v(231)
    and (n38, a[30], p[30]) ;   // shift.v(231)
    and (n39, a[31], p[31]) ;   // shift.v(231)
    not (n40, p[31]) ;   // shift.v(231)
    not (n41, p[30]) ;   // shift.v(231)
    not (n42, p[29]) ;   // shift.v(231)
    not (n43, p[28]) ;   // shift.v(231)
    not (n44, p[27]) ;   // shift.v(231)
    not (n45, p[26]) ;   // shift.v(231)
    not (n46, p[25]) ;   // shift.v(231)
    not (n47, p[24]) ;   // shift.v(231)
    not (n48, p[23]) ;   // shift.v(231)
    not (n49, p[22]) ;   // shift.v(231)
    not (n50, p[21]) ;   // shift.v(231)
    not (n51, p[20]) ;   // shift.v(231)
    not (n52, p[19]) ;   // shift.v(231)
    not (n53, p[18]) ;   // shift.v(231)
    not (n54, p[17]) ;   // shift.v(231)
    not (n55, p[16]) ;   // shift.v(231)
    not (n56, p[15]) ;   // shift.v(231)
    not (n57, p[14]) ;   // shift.v(231)
    not (n58, p[13]) ;   // shift.v(231)
    not (n59, p[12]) ;   // shift.v(231)
    not (n60, p[11]) ;   // shift.v(231)
    not (n61, p[10]) ;   // shift.v(231)
    not (n62, p[9]) ;   // shift.v(231)
    not (n63, p[8]) ;   // shift.v(231)
    not (n64, p[7]) ;   // shift.v(231)
    not (n65, p[6]) ;   // shift.v(231)
    not (n66, p[5]) ;   // shift.v(231)
    not (n67, p[4]) ;   // shift.v(231)
    not (n68, p[3]) ;   // shift.v(231)
    not (n69, p[2]) ;   // shift.v(231)
    not (n70, p[1]) ;   // shift.v(231)
    and (n71, s[30], n70) ;   // shift.v(231)
    and (n72, s[30], n69) ;   // shift.v(231)
    and (n73, s[30], n68) ;   // shift.v(231)
    and (n74, s[30], n67) ;   // shift.v(231)
    and (n75, s[30], n66) ;   // shift.v(231)
    and (n76, s[30], n65) ;   // shift.v(231)
    and (n77, s[30], n64) ;   // shift.v(231)
    and (n78, s[30], n63) ;   // shift.v(231)
    and (n79, s[30], n62) ;   // shift.v(231)
    and (n80, s[30], n61) ;   // shift.v(231)
    and (n81, s[30], n60) ;   // shift.v(231)
    and (n82, s[30], n59) ;   // shift.v(231)
    and (n83, s[30], n58) ;   // shift.v(231)
    and (n84, s[30], n57) ;   // shift.v(231)
    and (n85, s[30], n56) ;   // shift.v(231)
    and (n86, s[30], n55) ;   // shift.v(231)
    and (n87, s[30], n54) ;   // shift.v(231)
    and (n88, s[30], n53) ;   // shift.v(231)
    and (n89, s[30], n52) ;   // shift.v(231)
    and (n90, s[30], n51) ;   // shift.v(231)
    and (n91, s[30], n50) ;   // shift.v(231)
    and (n92, s[30], n49) ;   // shift.v(231)
    and (n93, s[30], n48) ;   // shift.v(231)
    and (n94, s[30], n47) ;   // shift.v(231)
    and (n95, s[30], n46) ;   // shift.v(231)
    and (n96, s[30], n45) ;   // shift.v(231)
    and (n97, s[30], n44) ;   // shift.v(231)
    and (n98, s[30], n43) ;   // shift.v(231)
    and (n99, s[30], n42) ;   // shift.v(231)
    and (n100, s[30], n41) ;   // shift.v(231)
    and (n101, s[30], n40) ;   // shift.v(231)
    or (q[1], n9, n71) ;   // shift.v(231)
    or (q[2], n10, n72) ;   // shift.v(231)
    or (q[3], n11, n73) ;   // shift.v(231)
    or (q[4], n12, n74) ;   // shift.v(231)
    or (q[5], n13, n75) ;   // shift.v(231)
    or (q[6], n14, n76) ;   // shift.v(231)
    or (q[7], n15, n77) ;   // shift.v(231)
    or (q[8], n16, n78) ;   // shift.v(231)
    or (q[9], n17, n79) ;   // shift.v(231)
    or (q[10], n18, n80) ;   // shift.v(231)
    or (q[11], n19, n81) ;   // shift.v(231)
    or (q[12], n20, n82) ;   // shift.v(231)
    or (q[13], n21, n83) ;   // shift.v(231)
    or (q[14], n22, n84) ;   // shift.v(231)
    or (q[15], n23, n85) ;   // shift.v(231)
    or (q[16], n24, n86) ;   // shift.v(231)
    or (q[17], n25, n87) ;   // shift.v(231)
    or (q[18], n26, n88) ;   // shift.v(231)
    or (q[19], n27, n89) ;   // shift.v(231)
    or (q[20], n28, n90) ;   // shift.v(231)
    or (q[21], n29, n91) ;   // shift.v(231)
    or (q[22], n30, n92) ;   // shift.v(231)
    or (q[23], n31, n93) ;   // shift.v(231)
    or (q[24], n32, n94) ;   // shift.v(231)
    or (q[25], n33, n95) ;   // shift.v(231)
    or (q[26], n34, n96) ;   // shift.v(231)
    or (q[27], n35, n97) ;   // shift.v(231)
    or (q[28], n36, n98) ;   // shift.v(231)
    or (q[29], n37, n99) ;   // shift.v(231)
    or (q[30], n38, n100) ;   // shift.v(231)
    or (q[31], n39, n101) ;   // shift.v(231)
    
endmodule

//
// Verific Verilog Description of module zmask_32
//

module zmask_32 (q, a, sla);   // shift.v(206)
    output [31:0]q;   // shift.v(210)
    input [31:0]a;   // shift.v(207)
    input sla;   // shift.v(208)
    
    
    or (q[0], sla, a[31]) ;   // shift.v(212)
    assign q[1] = sla ? a[31] : a[30];   // shift.v(216)
    assign q[2] = sla ? a[30] : a[29];   // shift.v(216)
    assign q[3] = sla ? a[29] : a[28];   // shift.v(216)
    assign q[4] = sla ? a[28] : a[27];   // shift.v(216)
    assign q[5] = sla ? a[27] : a[26];   // shift.v(216)
    assign q[6] = sla ? a[26] : a[25];   // shift.v(216)
    assign q[7] = sla ? a[25] : a[24];   // shift.v(216)
    assign q[8] = sla ? a[24] : a[23];   // shift.v(216)
    assign q[9] = sla ? a[23] : a[22];   // shift.v(216)
    assign q[10] = sla ? a[22] : a[21];   // shift.v(216)
    assign q[11] = sla ? a[21] : a[20];   // shift.v(216)
    assign q[12] = sla ? a[20] : a[19];   // shift.v(216)
    assign q[13] = sla ? a[19] : a[18];   // shift.v(216)
    assign q[14] = sla ? a[18] : a[17];   // shift.v(216)
    assign q[15] = sla ? a[17] : a[16];   // shift.v(216)
    assign q[16] = sla ? a[16] : a[15];   // shift.v(216)
    assign q[17] = sla ? a[15] : a[14];   // shift.v(216)
    assign q[18] = sla ? a[14] : a[13];   // shift.v(216)
    assign q[19] = sla ? a[13] : a[12];   // shift.v(216)
    assign q[20] = sla ? a[12] : a[11];   // shift.v(216)
    assign q[21] = sla ? a[11] : a[10];   // shift.v(216)
    assign q[22] = sla ? a[10] : a[9];   // shift.v(216)
    assign q[23] = sla ? a[9] : a[8];   // shift.v(216)
    assign q[24] = sla ? a[8] : a[7];   // shift.v(216)
    assign q[25] = sla ? a[7] : a[6];   // shift.v(216)
    assign q[26] = sla ? a[6] : a[5];   // shift.v(216)
    assign q[27] = sla ? a[5] : a[4];   // shift.v(216)
    assign q[28] = sla ? a[4] : a[3];   // shift.v(216)
    assign q[29] = sla ? a[3] : a[2];   // shift.v(216)
    assign q[30] = sla ? a[2] : a[1];   // shift.v(216)
    assign q[31] = sla ? a[1] : a[0];   // shift.v(216)
    
endmodule

//
// Verific Verilog Description of module ovf_32
//

module ovf_32 (q, a, f, sla);   // shift.v(192)
    output q;   // shift.v(197)
    input [31:0]a;   // shift.v(194)
    input [31:0]f;   // shift.v(193)
    input sla;   // shift.v(195)
    
    wire w1;   // shift.v(201)
    
    wire n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
        n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, 
        n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, 
        n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
        n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, 
        n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, 
        n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
        n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, 
        n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
        n95, n96;
    
    xor (n4, a[31], a[0]) ;   // shift.v(201)
    xor (n5, a[31], a[1]) ;   // shift.v(201)
    xor (n6, a[31], a[2]) ;   // shift.v(201)
    xor (n7, a[31], a[3]) ;   // shift.v(201)
    xor (n8, a[31], a[4]) ;   // shift.v(201)
    xor (n9, a[31], a[5]) ;   // shift.v(201)
    xor (n10, a[31], a[6]) ;   // shift.v(201)
    xor (n11, a[31], a[7]) ;   // shift.v(201)
    xor (n12, a[31], a[8]) ;   // shift.v(201)
    xor (n13, a[31], a[9]) ;   // shift.v(201)
    xor (n14, a[31], a[10]) ;   // shift.v(201)
    xor (n15, a[31], a[11]) ;   // shift.v(201)
    xor (n16, a[31], a[12]) ;   // shift.v(201)
    xor (n17, a[31], a[13]) ;   // shift.v(201)
    xor (n18, a[31], a[14]) ;   // shift.v(201)
    xor (n19, a[31], a[15]) ;   // shift.v(201)
    xor (n20, a[31], a[16]) ;   // shift.v(201)
    xor (n21, a[31], a[17]) ;   // shift.v(201)
    xor (n22, a[31], a[18]) ;   // shift.v(201)
    xor (n23, a[31], a[19]) ;   // shift.v(201)
    xor (n24, a[31], a[20]) ;   // shift.v(201)
    xor (n25, a[31], a[21]) ;   // shift.v(201)
    xor (n26, a[31], a[22]) ;   // shift.v(201)
    xor (n27, a[31], a[23]) ;   // shift.v(201)
    xor (n28, a[31], a[24]) ;   // shift.v(201)
    xor (n29, a[31], a[25]) ;   // shift.v(201)
    xor (n30, a[31], a[26]) ;   // shift.v(201)
    xor (n31, a[31], a[27]) ;   // shift.v(201)
    xor (n32, a[31], a[28]) ;   // shift.v(201)
    xor (n33, a[31], a[29]) ;   // shift.v(201)
    xor (n34, a[31], a[30]) ;   // shift.v(201)
    not (n35, f[31]) ;   // shift.v(201)
    not (n36, f[30]) ;   // shift.v(201)
    not (n37, f[29]) ;   // shift.v(201)
    not (n38, f[28]) ;   // shift.v(201)
    not (n39, f[27]) ;   // shift.v(201)
    not (n40, f[26]) ;   // shift.v(201)
    not (n41, f[25]) ;   // shift.v(201)
    not (n42, f[24]) ;   // shift.v(201)
    not (n43, f[23]) ;   // shift.v(201)
    not (n44, f[22]) ;   // shift.v(201)
    not (n45, f[21]) ;   // shift.v(201)
    not (n46, f[20]) ;   // shift.v(201)
    not (n47, f[19]) ;   // shift.v(201)
    not (n48, f[18]) ;   // shift.v(201)
    not (n49, f[17]) ;   // shift.v(201)
    not (n50, f[16]) ;   // shift.v(201)
    not (n51, f[15]) ;   // shift.v(201)
    not (n52, f[14]) ;   // shift.v(201)
    not (n53, f[13]) ;   // shift.v(201)
    not (n54, f[12]) ;   // shift.v(201)
    not (n55, f[11]) ;   // shift.v(201)
    not (n56, f[10]) ;   // shift.v(201)
    not (n57, f[9]) ;   // shift.v(201)
    not (n58, f[8]) ;   // shift.v(201)
    not (n59, f[7]) ;   // shift.v(201)
    not (n60, f[6]) ;   // shift.v(201)
    not (n61, f[5]) ;   // shift.v(201)
    not (n62, f[4]) ;   // shift.v(201)
    not (n63, f[3]) ;   // shift.v(201)
    not (n64, f[2]) ;   // shift.v(201)
    not (n65, f[1]) ;   // shift.v(201)
    and (n66, n4, n65) ;   // shift.v(201)
    and (n67, n5, n64) ;   // shift.v(201)
    and (n68, n6, n63) ;   // shift.v(201)
    and (n69, n7, n62) ;   // shift.v(201)
    and (n70, n8, n61) ;   // shift.v(201)
    and (n71, n9, n60) ;   // shift.v(201)
    and (n72, n10, n59) ;   // shift.v(201)
    and (n73, n11, n58) ;   // shift.v(201)
    and (n74, n12, n57) ;   // shift.v(201)
    and (n75, n13, n56) ;   // shift.v(201)
    and (n76, n14, n55) ;   // shift.v(201)
    and (n77, n15, n54) ;   // shift.v(201)
    and (n78, n16, n53) ;   // shift.v(201)
    and (n79, n17, n52) ;   // shift.v(201)
    and (n80, n18, n51) ;   // shift.v(201)
    and (n81, n19, n50) ;   // shift.v(201)
    and (n82, n20, n49) ;   // shift.v(201)
    and (n83, n21, n48) ;   // shift.v(201)
    and (n84, n22, n47) ;   // shift.v(201)
    and (n85, n23, n46) ;   // shift.v(201)
    and (n86, n24, n45) ;   // shift.v(201)
    and (n87, n25, n44) ;   // shift.v(201)
    and (n88, n26, n43) ;   // shift.v(201)
    and (n89, n27, n42) ;   // shift.v(201)
    and (n90, n28, n41) ;   // shift.v(201)
    and (n91, n29, n40) ;   // shift.v(201)
    and (n92, n30, n39) ;   // shift.v(201)
    and (n93, n31, n38) ;   // shift.v(201)
    and (n94, n32, n37) ;   // shift.v(201)
    and (n95, n33, n36) ;   // shift.v(201)
    and (n96, n34, n35) ;   // shift.v(201)
    or (w1, n96, n95, n94, n93, n92, n91, n90, n89, n88, 
        n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69, n68, 
        n67, n66) ;   // shift.v(201)
    and (q, sla, w1) ;   // shift.v(203)
    
endmodule

//
// Verific Verilog Description of module mul_32
//

module mul_32 (q1, q2, ov, z, a, b);   // alu.v(23)
    output [31:0]q1;   // alu.v(26)
    output [31:0]q2;   // alu.v(26)
    output ov;   // alu.v(27)
    output z;   // alu.v(27)
    input [31:0]a;   // alu.v(24)
    input [31:0]b;   // alu.v(24)
    
    
    mult_32 m0 (.a({a}), .b({b}), .m({q2, q1}));   // alu.v(33)
    or (ov, q2[31], q2[30], q2[29], q2[28], q2[27], q2[26], q2[25], 
            q2[24], q2[23], q2[22], q2[21], q2[20], q2[19], q2[18], 
            q2[17], q2[16], q2[15], q2[14], q2[13], q2[12], q2[11], 
            q2[10], q2[9], q2[8], q2[7], q2[6], q2[5], q2[4], 
            q2[3], q2[2], q2[1], q2[0]) ;   // alu.v(35)
    nor (z, q2[31], q2[30], q2[29], q2[28], q2[27], q2[26], q2[25], 
            q2[24], q2[23], q2[22], q2[21], q2[20], q2[19], q2[18], 
            q2[17], q2[16], q2[15], q2[14], q2[13], q2[12], q2[11], 
            q2[10], q2[9], q2[8], q2[7], q2[6], q2[5], q2[4], 
            q2[3], q2[2], q2[1], q2[0], q1[31], q1[30], q1[29], 
            q1[28], q1[27], q1[26], q1[25], q1[24], q1[23], q1[22], 
            q1[21], q1[20], q1[19], q1[18], q1[17], q1[16], q1[15], 
            q1[14], q1[13], q1[12], q1[11], q1[10], q1[9], q1[8], 
            q1[7], q1[6], q1[5], q1[4], q1[3], q1[2], q1[1], q1[0]) ;   // alu.v(36)
    
endmodule

//
// Verific Verilog Description of module mult_32
//

module mult_32 (a, b, m);   // mult.v(36)
    input [31:0]a;   // mult.v(37)
    input [31:0]b;   // mult.v(38)
    output [63:0]m;   // mult.v(40)
    
    wire wand_28;   // mult.v(43)
    wire wand_59;   // mult.v(44)
    wire wha_s_0;   // mult.v(45)
    wire wha_c_0;   // mult.v(45)
    wire wand_29;   // mult.v(46)
    wire wand_60;   // mult.v(47)
    wire wand_91;   // mult.v(48)
    wire wfa_s_0;   // mult.v(49)
    wire wfa_cout_0;   // mult.v(49)
    wire wand_122;   // mult.v(50)
    wire wand_153;   // mult.v(51)
    wire wha_s_1;   // mult.v(52)
    wire wha_c_1;   // mult.v(52)
    wire wand_30;   // mult.v(53)
    wire wand_61;   // mult.v(54)
    wire wand_92;   // mult.v(55)
    wire wfa_s_1;   // mult.v(56)
    wire wfa_cout_1;   // mult.v(56)
    wire wand_123;   // mult.v(57)
    wire wand_154;   // mult.v(58)
    wire wand_185;   // mult.v(59)
    wire wfa_s_2;   // mult.v(60)
    wire wfa_cout_2;   // mult.v(60)
    wire wand_216;   // mult.v(61)
    wire wand_247;   // mult.v(62)
    wire wha_s_2;   // mult.v(63)
    wire wha_c_2;   // mult.v(63)
    wire wand_31;   // mult.v(64)
    wire wand_62;   // mult.v(65)
    wire wand_93;   // mult.v(66)
    wire wfa_s_3;   // mult.v(67)
    wire wfa_cout_3;   // mult.v(67)
    wire wand_124;   // mult.v(68)
    wire wand_155;   // mult.v(69)
    wire wand_186;   // mult.v(70)
    wire wfa_s_4;   // mult.v(71)
    wire wfa_cout_4;   // mult.v(71)
    wire wand_217;   // mult.v(72)
    wire wand_248;   // mult.v(73)
    wire wand_279;   // mult.v(74)
    wire wfa_s_5;   // mult.v(75)
    wire wfa_cout_5;   // mult.v(75)
    wire wand_310;   // mult.v(76)
    wire wand_341;   // mult.v(77)
    wire wha_s_3;   // mult.v(78)
    wire wha_c_3;   // mult.v(78)
    wire wand_63;   // mult.v(79)
    wire wand_94;   // mult.v(80)
    wire wand_125;   // mult.v(81)
    wire wfa_s_6;   // mult.v(82)
    wire wfa_cout_6;   // mult.v(82)
    wire wand_156;   // mult.v(83)
    wire wand_187;   // mult.v(84)
    wire wand_218;   // mult.v(85)
    wire wfa_s_7;   // mult.v(86)
    wire wfa_cout_7;   // mult.v(86)
    wire wand_249;   // mult.v(87)
    wire wand_280;   // mult.v(88)
    wire wand_311;   // mult.v(89)
    wire wfa_s_8;   // mult.v(90)
    wire wfa_cout_8;   // mult.v(90)
    wire wand_342;   // mult.v(91)
    wire wand_373;   // mult.v(92)
    wire wha_s_4;   // mult.v(93)
    wire wha_c_4;   // mult.v(93)
    wire wand_95;   // mult.v(94)
    wire wand_126;   // mult.v(95)
    wire wand_157;   // mult.v(96)
    wire wfa_s_9;   // mult.v(97)
    wire wfa_cout_9;   // mult.v(97)
    wire wand_188;   // mult.v(98)
    wire wand_219;   // mult.v(99)
    wire wand_250;   // mult.v(100)
    wire wfa_s_10;   // mult.v(101)
    wire wfa_cout_10;   // mult.v(101)
    wire wand_281;   // mult.v(102)
    wire wand_312;   // mult.v(103)
    wire wand_343;   // mult.v(104)
    wire wfa_s_11;   // mult.v(105)
    wire wfa_cout_11;   // mult.v(105)
    wire wand_127;   // mult.v(106)
    wire wand_158;   // mult.v(107)
    wire wand_189;   // mult.v(108)
    wire wfa_s_12;   // mult.v(109)
    wire wfa_cout_12;   // mult.v(109)
    wire wand_220;   // mult.v(110)
    wire wand_251;   // mult.v(111)
    wire wand_282;   // mult.v(112)
    wire wfa_s_13;   // mult.v(113)
    wire wfa_cout_13;   // mult.v(113)
    wire wand_159;   // mult.v(114)
    wire wand_190;   // mult.v(115)
    wire wand_221;   // mult.v(116)
    wire wfa_s_14;   // mult.v(117)
    wire wfa_cout_14;   // mult.v(117)
    wire wand_19;   // mult.v(118)
    wire wand_50;   // mult.v(119)
    wire wha_s_5;   // mult.v(120)
    wire wha_c_5;   // mult.v(120)
    wire wand_20;   // mult.v(121)
    wire wand_51;   // mult.v(122)
    wire wand_82;   // mult.v(123)
    wire wfa_s_15;   // mult.v(124)
    wire wfa_cout_15;   // mult.v(124)
    wire wand_113;   // mult.v(125)
    wire wand_144;   // mult.v(126)
    wire wha_s_6;   // mult.v(127)
    wire wha_c_6;   // mult.v(127)
    wire wand_21;   // mult.v(128)
    wire wand_52;   // mult.v(129)
    wire wand_83;   // mult.v(130)
    wire wfa_s_16;   // mult.v(131)
    wire wfa_cout_16;   // mult.v(131)
    wire wand_114;   // mult.v(132)
    wire wand_145;   // mult.v(133)
    wire wand_176;   // mult.v(134)
    wire wfa_s_17;   // mult.v(135)
    wire wfa_cout_17;   // mult.v(135)
    wire wand_207;   // mult.v(136)
    wire wand_238;   // mult.v(137)
    wire wha_s_7;   // mult.v(138)
    wire wha_c_7;   // mult.v(138)
    wire wand_22;   // mult.v(139)
    wire wand_53;   // mult.v(140)
    wire wand_84;   // mult.v(141)
    wire wfa_s_18;   // mult.v(142)
    wire wfa_cout_18;   // mult.v(142)
    wire wand_115;   // mult.v(143)
    wire wand_146;   // mult.v(144)
    wire wand_177;   // mult.v(145)
    wire wfa_s_19;   // mult.v(146)
    wire wfa_cout_19;   // mult.v(146)
    wire wand_208;   // mult.v(147)
    wire wand_239;   // mult.v(148)
    wire wand_270;   // mult.v(149)
    wire wfa_s_20;   // mult.v(150)
    wire wfa_cout_20;   // mult.v(150)
    wire wand_301;   // mult.v(151)
    wire wand_332;   // mult.v(152)
    wire wha_s_8;   // mult.v(153)
    wire wha_c_8;   // mult.v(153)
    wire wand_23;   // mult.v(154)
    wire wand_54;   // mult.v(155)
    wire wand_85;   // mult.v(156)
    wire wfa_s_21;   // mult.v(157)
    wire wfa_cout_21;   // mult.v(157)
    wire wand_116;   // mult.v(158)
    wire wand_147;   // mult.v(159)
    wire wand_178;   // mult.v(160)
    wire wfa_s_22;   // mult.v(161)
    wire wfa_cout_22;   // mult.v(161)
    wire wand_209;   // mult.v(162)
    wire wand_240;   // mult.v(163)
    wire wand_271;   // mult.v(164)
    wire wfa_s_23;   // mult.v(165)
    wire wfa_cout_23;   // mult.v(165)
    wire wand_302;   // mult.v(166)
    wire wand_333;   // mult.v(167)
    wire wand_364;   // mult.v(168)
    wire wfa_s_24;   // mult.v(169)
    wire wfa_cout_24;   // mult.v(169)
    wire wand_395;   // mult.v(170)
    wire wand_426;   // mult.v(171)
    wire wha_s_9;   // mult.v(172)
    wire wha_c_9;   // mult.v(172)
    wire wand_24;   // mult.v(173)
    wire wand_55;   // mult.v(174)
    wire wand_86;   // mult.v(175)
    wire wfa_s_25;   // mult.v(176)
    wire wfa_cout_25;   // mult.v(176)
    wire wand_117;   // mult.v(177)
    wire wand_148;   // mult.v(178)
    wire wand_179;   // mult.v(179)
    wire wfa_s_26;   // mult.v(180)
    wire wfa_cout_26;   // mult.v(180)
    wire wand_210;   // mult.v(181)
    wire wand_241;   // mult.v(182)
    wire wand_272;   // mult.v(183)
    wire wfa_s_27;   // mult.v(184)
    wire wfa_cout_27;   // mult.v(184)
    wire wand_303;   // mult.v(185)
    wire wand_334;   // mult.v(186)
    wire wand_365;   // mult.v(187)
    wire wfa_s_28;   // mult.v(188)
    wire wfa_cout_28;   // mult.v(188)
    wire wand_396;   // mult.v(189)
    wire wand_427;   // mult.v(190)
    wire wand_458;   // mult.v(191)
    wire wfa_s_29;   // mult.v(192)
    wire wfa_cout_29;   // mult.v(192)
    wire wand_489;   // mult.v(193)
    wire wand_520;   // mult.v(194)
    wire wha_s_10;   // mult.v(195)
    wire wha_c_10;   // mult.v(195)
    wire wand_25;   // mult.v(196)
    wire wand_56;   // mult.v(197)
    wire wand_87;   // mult.v(198)
    wire wfa_s_30;   // mult.v(199)
    wire wfa_cout_30;   // mult.v(199)
    wire wand_118;   // mult.v(200)
    wire wand_149;   // mult.v(201)
    wire wand_180;   // mult.v(202)
    wire wfa_s_31;   // mult.v(203)
    wire wfa_cout_31;   // mult.v(203)
    wire wand_211;   // mult.v(204)
    wire wand_242;   // mult.v(205)
    wire wand_273;   // mult.v(206)
    wire wfa_s_32;   // mult.v(207)
    wire wfa_cout_32;   // mult.v(207)
    wire wand_304;   // mult.v(208)
    wire wand_335;   // mult.v(209)
    wire wand_366;   // mult.v(210)
    wire wfa_s_33;   // mult.v(211)
    wire wfa_cout_33;   // mult.v(211)
    wire wand_397;   // mult.v(212)
    wire wand_428;   // mult.v(213)
    wire wand_459;   // mult.v(214)
    wire wfa_s_34;   // mult.v(215)
    wire wfa_cout_34;   // mult.v(215)
    wire wand_490;   // mult.v(216)
    wire wand_521;   // mult.v(217)
    wire wand_552;   // mult.v(218)
    wire wfa_s_35;   // mult.v(219)
    wire wfa_cout_35;   // mult.v(219)
    wire wand_583;   // mult.v(220)
    wire wand_614;   // mult.v(221)
    wire wha_s_11;   // mult.v(222)
    wire wha_c_11;   // mult.v(222)
    wire wand_26;   // mult.v(223)
    wire wand_57;   // mult.v(224)
    wire wand_88;   // mult.v(225)
    wire wfa_s_36;   // mult.v(226)
    wire wfa_cout_36;   // mult.v(226)
    wire wand_119;   // mult.v(227)
    wire wand_150;   // mult.v(228)
    wire wand_181;   // mult.v(229)
    wire wfa_s_37;   // mult.v(230)
    wire wfa_cout_37;   // mult.v(230)
    wire wand_212;   // mult.v(231)
    wire wand_243;   // mult.v(232)
    wire wand_274;   // mult.v(233)
    wire wfa_s_38;   // mult.v(234)
    wire wfa_cout_38;   // mult.v(234)
    wire wand_305;   // mult.v(235)
    wire wand_336;   // mult.v(236)
    wire wand_367;   // mult.v(237)
    wire wfa_s_39;   // mult.v(238)
    wire wfa_cout_39;   // mult.v(238)
    wire wand_398;   // mult.v(239)
    wire wand_429;   // mult.v(240)
    wire wand_460;   // mult.v(241)
    wire wfa_s_40;   // mult.v(242)
    wire wfa_cout_40;   // mult.v(242)
    wire wand_491;   // mult.v(243)
    wire wand_522;   // mult.v(244)
    wire wand_553;   // mult.v(245)
    wire wfa_s_41;   // mult.v(246)
    wire wfa_cout_41;   // mult.v(246)
    wire wand_584;   // mult.v(247)
    wire wand_615;   // mult.v(248)
    wire wand_646;   // mult.v(249)
    wire wfa_s_42;   // mult.v(250)
    wire wfa_cout_42;   // mult.v(250)
    wire wand_677;   // mult.v(251)
    wire wand_708;   // mult.v(252)
    wire wha_s_12;   // mult.v(253)
    wire wha_c_12;   // mult.v(253)
    wire wand_27;   // mult.v(254)
    wire wand_58;   // mult.v(255)
    wire wand_89;   // mult.v(256)
    wire wfa_s_43;   // mult.v(257)
    wire wfa_cout_43;   // mult.v(257)
    wire wand_120;   // mult.v(258)
    wire wand_151;   // mult.v(259)
    wire wand_182;   // mult.v(260)
    wire wfa_s_44;   // mult.v(261)
    wire wfa_cout_44;   // mult.v(261)
    wire wand_213;   // mult.v(262)
    wire wand_244;   // mult.v(263)
    wire wand_275;   // mult.v(264)
    wire wfa_s_45;   // mult.v(265)
    wire wfa_cout_45;   // mult.v(265)
    wire wand_306;   // mult.v(266)
    wire wand_337;   // mult.v(267)
    wire wand_368;   // mult.v(268)
    wire wfa_s_46;   // mult.v(269)
    wire wfa_cout_46;   // mult.v(269)
    wire wand_399;   // mult.v(270)
    wire wand_430;   // mult.v(271)
    wire wand_461;   // mult.v(272)
    wire wfa_s_47;   // mult.v(273)
    wire wfa_cout_47;   // mult.v(273)
    wire wand_492;   // mult.v(274)
    wire wand_523;   // mult.v(275)
    wire wand_554;   // mult.v(276)
    wire wfa_s_48;   // mult.v(277)
    wire wfa_cout_48;   // mult.v(277)
    wire wand_585;   // mult.v(278)
    wire wand_616;   // mult.v(279)
    wire wand_647;   // mult.v(280)
    wire wfa_s_49;   // mult.v(281)
    wire wfa_cout_49;   // mult.v(281)
    wire wand_678;   // mult.v(282)
    wire wand_709;   // mult.v(283)
    wire wand_740;   // mult.v(284)
    wire wfa_s_50;   // mult.v(285)
    wire wfa_cout_50;   // mult.v(285)
    wire wand_771;   // mult.v(286)
    wire wand_802;   // mult.v(287)
    wire wha_s_13;   // mult.v(288)
    wire wha_c_13;   // mult.v(288)
    wire wand_90;   // mult.v(289)
    wire wand_121;   // mult.v(290)
    wire wand_152;   // mult.v(291)
    wire wfa_s_51;   // mult.v(292)
    wire wfa_cout_51;   // mult.v(292)
    wire wand_183;   // mult.v(293)
    wire wand_214;   // mult.v(294)
    wire wand_245;   // mult.v(295)
    wire wfa_s_52;   // mult.v(296)
    wire wfa_cout_52;   // mult.v(296)
    wire wand_276;   // mult.v(297)
    wire wand_307;   // mult.v(298)
    wire wand_338;   // mult.v(299)
    wire wfa_s_53;   // mult.v(300)
    wire wfa_cout_53;   // mult.v(300)
    wire wand_369;   // mult.v(301)
    wire wand_400;   // mult.v(302)
    wire wand_431;   // mult.v(303)
    wire wfa_s_54;   // mult.v(304)
    wire wfa_cout_54;   // mult.v(304)
    wire wand_462;   // mult.v(305)
    wire wand_493;   // mult.v(306)
    wire wand_524;   // mult.v(307)
    wire wfa_s_55;   // mult.v(308)
    wire wfa_cout_55;   // mult.v(308)
    wire wand_555;   // mult.v(309)
    wire wand_586;   // mult.v(310)
    wire wand_617;   // mult.v(311)
    wire wfa_s_56;   // mult.v(312)
    wire wfa_cout_56;   // mult.v(312)
    wire wand_648;   // mult.v(313)
    wire wand_679;   // mult.v(314)
    wire wand_710;   // mult.v(315)
    wire wfa_s_57;   // mult.v(316)
    wire wfa_cout_57;   // mult.v(316)
    wire wand_741;   // mult.v(317)
    wire wand_772;   // mult.v(318)
    wire wand_803;   // mult.v(319)
    wire wfa_s_58;   // mult.v(320)
    wire wfa_cout_58;   // mult.v(320)
    wire wand_834;   // mult.v(321)
    wire wand_865;   // mult.v(322)
    wire wand_896;   // mult.v(323)
    wire wfa_s_59;   // mult.v(324)
    wire wfa_cout_59;   // mult.v(324)
    wire wand_184;   // mult.v(325)
    wire wand_215;   // mult.v(326)
    wire wand_246;   // mult.v(327)
    wire wfa_s_60;   // mult.v(328)
    wire wfa_cout_60;   // mult.v(328)
    wire wand_277;   // mult.v(329)
    wire wand_308;   // mult.v(330)
    wire wand_339;   // mult.v(331)
    wire wfa_s_61;   // mult.v(332)
    wire wfa_cout_61;   // mult.v(332)
    wire wand_370;   // mult.v(333)
    wire wand_401;   // mult.v(334)
    wire wand_432;   // mult.v(335)
    wire wfa_s_62;   // mult.v(336)
    wire wfa_cout_62;   // mult.v(336)
    wire wand_463;   // mult.v(337)
    wire wand_494;   // mult.v(338)
    wire wand_525;   // mult.v(339)
    wire wfa_s_63;   // mult.v(340)
    wire wfa_cout_63;   // mult.v(340)
    wire wand_556;   // mult.v(341)
    wire wand_587;   // mult.v(342)
    wire wand_618;   // mult.v(343)
    wire wfa_s_64;   // mult.v(344)
    wire wfa_cout_64;   // mult.v(344)
    wire wand_649;   // mult.v(345)
    wire wand_680;   // mult.v(346)
    wire wand_711;   // mult.v(347)
    wire wfa_s_65;   // mult.v(348)
    wire wfa_cout_65;   // mult.v(348)
    wire wand_742;   // mult.v(349)
    wire wand_773;   // mult.v(350)
    wire wand_804;   // mult.v(351)
    wire wfa_s_66;   // mult.v(352)
    wire wfa_cout_66;   // mult.v(352)
    wire wand_835;   // mult.v(353)
    wire wand_866;   // mult.v(354)
    wire wand_897;   // mult.v(355)
    wire wfa_s_67;   // mult.v(356)
    wire wfa_cout_67;   // mult.v(356)
    wire wand_928;   // mult.v(357)
    wire wfa_s_68;   // mult.v(358)
    wire wfa_cout_68;   // mult.v(358)
    wire wand_278;   // mult.v(359)
    wire wand_309;   // mult.v(360)
    wire wand_340;   // mult.v(361)
    wire wfa_s_69;   // mult.v(362)
    wire wfa_cout_69;   // mult.v(362)
    wire wand_371;   // mult.v(363)
    wire wand_402;   // mult.v(364)
    wire wand_433;   // mult.v(365)
    wire wfa_s_70;   // mult.v(366)
    wire wfa_cout_70;   // mult.v(366)
    wire wand_464;   // mult.v(367)
    wire wand_495;   // mult.v(368)
    wire wand_526;   // mult.v(369)
    wire wfa_s_71;   // mult.v(370)
    wire wfa_cout_71;   // mult.v(370)
    wire wand_557;   // mult.v(371)
    wire wand_588;   // mult.v(372)
    wire wand_619;   // mult.v(373)
    wire wfa_s_72;   // mult.v(374)
    wire wfa_cout_72;   // mult.v(374)
    wire wand_650;   // mult.v(375)
    wire wand_681;   // mult.v(376)
    wire wand_712;   // mult.v(377)
    wire wfa_s_73;   // mult.v(378)
    wire wfa_cout_73;   // mult.v(378)
    wire wand_743;   // mult.v(379)
    wire wand_774;   // mult.v(380)
    wire wand_805;   // mult.v(381)
    wire wfa_s_74;   // mult.v(382)
    wire wfa_cout_74;   // mult.v(382)
    wire wand_836;   // mult.v(383)
    wire wand_867;   // mult.v(384)
    wire wand_898;   // mult.v(385)
    wire wfa_s_75;   // mult.v(386)
    wire wfa_cout_75;   // mult.v(386)
    wire wand_929;   // mult.v(387)
    wire wand_960;   // mult.v(388)
    wire wfa_s_76;   // mult.v(389)
    wire wfa_cout_76;   // mult.v(389)
    wire wfa_s_77;   // mult.v(390)
    wire wfa_cout_77;   // mult.v(390)
    wire wand_372;   // mult.v(391)
    wire wand_403;   // mult.v(392)
    wire wand_434;   // mult.v(393)
    wire wfa_s_78;   // mult.v(394)
    wire wfa_cout_78;   // mult.v(394)
    wire wand_465;   // mult.v(395)
    wire wand_496;   // mult.v(396)
    wire wand_527;   // mult.v(397)
    wire wfa_s_79;   // mult.v(398)
    wire wfa_cout_79;   // mult.v(398)
    wire wand_558;   // mult.v(399)
    wire wand_589;   // mult.v(400)
    wire wand_620;   // mult.v(401)
    wire wfa_s_80;   // mult.v(402)
    wire wfa_cout_80;   // mult.v(402)
    wire wand_651;   // mult.v(403)
    wire wand_682;   // mult.v(404)
    wire wand_713;   // mult.v(405)
    wire wfa_s_81;   // mult.v(406)
    wire wfa_cout_81;   // mult.v(406)
    wire wand_744;   // mult.v(407)
    wire wand_775;   // mult.v(408)
    wire wand_806;   // mult.v(409)
    wire wfa_s_82;   // mult.v(410)
    wire wfa_cout_82;   // mult.v(410)
    wire wand_837;   // mult.v(411)
    wire wand_868;   // mult.v(412)
    wire wand_899;   // mult.v(413)
    wire wfa_s_83;   // mult.v(414)
    wire wfa_cout_83;   // mult.v(414)
    wire wand_930;   // mult.v(415)
    wire wand_961;   // mult.v(416)
    wire wand_992;   // mult.v(417)
    wire wfa_s_84;   // mult.v(418)
    wire wfa_cout_84;   // mult.v(418)
    wire wfa_s_85;   // mult.v(419)
    wire wfa_cout_85;   // mult.v(419)
    wire wfa_s_86;   // mult.v(420)
    wire wfa_cout_86;   // mult.v(420)
    wire wand_404;   // mult.v(421)
    wire wand_435;   // mult.v(422)
    wire wand_466;   // mult.v(423)
    wire wfa_s_87;   // mult.v(424)
    wire wfa_cout_87;   // mult.v(424)
    wire wand_497;   // mult.v(425)
    wire wand_528;   // mult.v(426)
    wire wand_559;   // mult.v(427)
    wire wfa_s_88;   // mult.v(428)
    wire wfa_cout_88;   // mult.v(428)
    wire wand_590;   // mult.v(429)
    wire wand_621;   // mult.v(430)
    wire wand_652;   // mult.v(431)
    wire wfa_s_89;   // mult.v(432)
    wire wfa_cout_89;   // mult.v(432)
    wire wand_683;   // mult.v(433)
    wire wand_714;   // mult.v(434)
    wire wand_745;   // mult.v(435)
    wire wfa_s_90;   // mult.v(436)
    wire wfa_cout_90;   // mult.v(436)
    wire wand_776;   // mult.v(437)
    wire wand_807;   // mult.v(438)
    wire wand_838;   // mult.v(439)
    wire wfa_s_91;   // mult.v(440)
    wire wfa_cout_91;   // mult.v(440)
    wire wand_869;   // mult.v(441)
    wire wand_900;   // mult.v(442)
    wire wand_931;   // mult.v(443)
    wire wfa_s_92;   // mult.v(444)
    wire wfa_cout_92;   // mult.v(444)
    wire wand_962;   // mult.v(445)
    wire wand_993;   // mult.v(446)
    wire wfa_s_93;   // mult.v(447)
    wire wfa_cout_93;   // mult.v(447)
    wire wfa_s_94;   // mult.v(448)
    wire wfa_cout_94;   // mult.v(448)
    wire wfa_s_95;   // mult.v(449)
    wire wfa_cout_95;   // mult.v(449)
    wire wand_374;   // mult.v(450)
    wire wand_405;   // mult.v(451)
    wire wand_436;   // mult.v(452)
    wire wfa_s_96;   // mult.v(453)
    wire wfa_cout_96;   // mult.v(453)
    wire wand_467;   // mult.v(454)
    wire wand_498;   // mult.v(455)
    wire wand_529;   // mult.v(456)
    wire wfa_s_97;   // mult.v(457)
    wire wfa_cout_97;   // mult.v(457)
    wire wand_560;   // mult.v(458)
    wire wand_591;   // mult.v(459)
    wire wand_622;   // mult.v(460)
    wire wfa_s_98;   // mult.v(461)
    wire wfa_cout_98;   // mult.v(461)
    wire wand_653;   // mult.v(462)
    wire wand_684;   // mult.v(463)
    wire wand_715;   // mult.v(464)
    wire wfa_s_99;   // mult.v(465)
    wire wfa_cout_99;   // mult.v(465)
    wire wand_746;   // mult.v(466)
    wire wand_777;   // mult.v(467)
    wire wand_808;   // mult.v(468)
    wire wfa_s_100;   // mult.v(469)
    wire wfa_cout_100;   // mult.v(469)
    wire wand_839;   // mult.v(470)
    wire wand_870;   // mult.v(471)
    wire wand_901;   // mult.v(472)
    wire wfa_s_101;   // mult.v(473)
    wire wfa_cout_101;   // mult.v(473)
    wire wand_932;   // mult.v(474)
    wire wand_963;   // mult.v(475)
    wire wand_994;   // mult.v(476)
    wire wfa_s_102;   // mult.v(477)
    wire wfa_cout_102;   // mult.v(477)
    wire wfa_s_103;   // mult.v(478)
    wire wfa_cout_103;   // mult.v(478)
    wire wfa_s_104;   // mult.v(479)
    wire wfa_cout_104;   // mult.v(479)
    wire wand_313;   // mult.v(480)
    wire wand_344;   // mult.v(481)
    wire wand_375;   // mult.v(482)
    wire wfa_s_105;   // mult.v(483)
    wire wfa_cout_105;   // mult.v(483)
    wire wand_406;   // mult.v(484)
    wire wand_437;   // mult.v(485)
    wire wand_468;   // mult.v(486)
    wire wfa_s_106;   // mult.v(487)
    wire wfa_cout_106;   // mult.v(487)
    wire wand_499;   // mult.v(488)
    wire wand_530;   // mult.v(489)
    wire wand_561;   // mult.v(490)
    wire wfa_s_107;   // mult.v(491)
    wire wfa_cout_107;   // mult.v(491)
    wire wand_592;   // mult.v(492)
    wire wand_623;   // mult.v(493)
    wire wand_654;   // mult.v(494)
    wire wfa_s_108;   // mult.v(495)
    wire wfa_cout_108;   // mult.v(495)
    wire wand_685;   // mult.v(496)
    wire wand_716;   // mult.v(497)
    wire wand_747;   // mult.v(498)
    wire wfa_s_109;   // mult.v(499)
    wire wfa_cout_109;   // mult.v(499)
    wire wand_778;   // mult.v(500)
    wire wand_809;   // mult.v(501)
    wire wand_840;   // mult.v(502)
    wire wfa_s_110;   // mult.v(503)
    wire wfa_cout_110;   // mult.v(503)
    wire wand_871;   // mult.v(504)
    wire wand_902;   // mult.v(505)
    wire wand_933;   // mult.v(506)
    wire wfa_s_111;   // mult.v(507)
    wire wfa_cout_111;   // mult.v(507)
    wire wand_964;   // mult.v(508)
    wire wand_995;   // mult.v(509)
    wire wfa_s_112;   // mult.v(510)
    wire wfa_cout_112;   // mult.v(510)
    wire wfa_s_113;   // mult.v(511)
    wire wfa_cout_113;   // mult.v(511)
    wire wand_252;   // mult.v(512)
    wire wand_283;   // mult.v(513)
    wire wand_314;   // mult.v(514)
    wire wfa_s_114;   // mult.v(515)
    wire wfa_cout_114;   // mult.v(515)
    wire wand_345;   // mult.v(516)
    wire wand_376;   // mult.v(517)
    wire wand_407;   // mult.v(518)
    wire wfa_s_115;   // mult.v(519)
    wire wfa_cout_115;   // mult.v(519)
    wire wand_438;   // mult.v(520)
    wire wand_469;   // mult.v(521)
    wire wand_500;   // mult.v(522)
    wire wfa_s_116;   // mult.v(523)
    wire wfa_cout_116;   // mult.v(523)
    wire wand_531;   // mult.v(524)
    wire wand_562;   // mult.v(525)
    wire wand_593;   // mult.v(526)
    wire wfa_s_117;   // mult.v(527)
    wire wfa_cout_117;   // mult.v(527)
    wire wand_624;   // mult.v(528)
    wire wand_655;   // mult.v(529)
    wire wand_686;   // mult.v(530)
    wire wfa_s_118;   // mult.v(531)
    wire wfa_cout_118;   // mult.v(531)
    wire wand_717;   // mult.v(532)
    wire wand_748;   // mult.v(533)
    wire wand_779;   // mult.v(534)
    wire wfa_s_119;   // mult.v(535)
    wire wfa_cout_119;   // mult.v(535)
    wire wand_810;   // mult.v(536)
    wire wand_841;   // mult.v(537)
    wire wand_872;   // mult.v(538)
    wire wfa_s_120;   // mult.v(539)
    wire wfa_cout_120;   // mult.v(539)
    wire wand_903;   // mult.v(540)
    wire wand_934;   // mult.v(541)
    wire wand_965;   // mult.v(542)
    wire wfa_s_121;   // mult.v(543)
    wire wfa_cout_121;   // mult.v(543)
    wire wand_996;   // mult.v(544)
    wire wfa_s_122;   // mult.v(545)
    wire wfa_cout_122;   // mult.v(545)
    wire wand_191;   // mult.v(546)
    wire wand_222;   // mult.v(547)
    wire wand_253;   // mult.v(548)
    wire wfa_s_123;   // mult.v(549)
    wire wfa_cout_123;   // mult.v(549)
    wire wand_284;   // mult.v(550)
    wire wand_315;   // mult.v(551)
    wire wand_346;   // mult.v(552)
    wire wfa_s_124;   // mult.v(553)
    wire wfa_cout_124;   // mult.v(553)
    wire wand_377;   // mult.v(554)
    wire wand_408;   // mult.v(555)
    wire wand_439;   // mult.v(556)
    wire wfa_s_125;   // mult.v(557)
    wire wfa_cout_125;   // mult.v(557)
    wire wand_470;   // mult.v(558)
    wire wand_501;   // mult.v(559)
    wire wand_532;   // mult.v(560)
    wire wfa_s_126;   // mult.v(561)
    wire wfa_cout_126;   // mult.v(561)
    wire wand_563;   // mult.v(562)
    wire wand_594;   // mult.v(563)
    wire wand_625;   // mult.v(564)
    wire wfa_s_127;   // mult.v(565)
    wire wfa_cout_127;   // mult.v(565)
    wire wand_656;   // mult.v(566)
    wire wand_687;   // mult.v(567)
    wire wand_718;   // mult.v(568)
    wire wfa_s_128;   // mult.v(569)
    wire wfa_cout_128;   // mult.v(569)
    wire wand_749;   // mult.v(570)
    wire wand_780;   // mult.v(571)
    wire wand_811;   // mult.v(572)
    wire wfa_s_129;   // mult.v(573)
    wire wfa_cout_129;   // mult.v(573)
    wire wand_842;   // mult.v(574)
    wire wand_873;   // mult.v(575)
    wire wand_904;   // mult.v(576)
    wire wfa_s_130;   // mult.v(577)
    wire wfa_cout_130;   // mult.v(577)
    wire wand_935;   // mult.v(578)
    wire wand_966;   // mult.v(579)
    wire wand_997;   // mult.v(580)
    wire wfa_s_131;   // mult.v(581)
    wire wfa_cout_131;   // mult.v(581)
    wire wand_223;   // mult.v(582)
    wire wand_254;   // mult.v(583)
    wire wand_285;   // mult.v(584)
    wire wfa_s_132;   // mult.v(585)
    wire wfa_cout_132;   // mult.v(585)
    wire wand_316;   // mult.v(586)
    wire wand_347;   // mult.v(587)
    wire wand_378;   // mult.v(588)
    wire wfa_s_133;   // mult.v(589)
    wire wfa_cout_133;   // mult.v(589)
    wire wand_409;   // mult.v(590)
    wire wand_440;   // mult.v(591)
    wire wand_471;   // mult.v(592)
    wire wfa_s_134;   // mult.v(593)
    wire wfa_cout_134;   // mult.v(593)
    wire wand_502;   // mult.v(594)
    wire wand_533;   // mult.v(595)
    wire wand_564;   // mult.v(596)
    wire wfa_s_135;   // mult.v(597)
    wire wfa_cout_135;   // mult.v(597)
    wire wand_595;   // mult.v(598)
    wire wand_626;   // mult.v(599)
    wire wand_657;   // mult.v(600)
    wire wfa_s_136;   // mult.v(601)
    wire wfa_cout_136;   // mult.v(601)
    wire wand_688;   // mult.v(602)
    wire wand_719;   // mult.v(603)
    wire wand_750;   // mult.v(604)
    wire wfa_s_137;   // mult.v(605)
    wire wfa_cout_137;   // mult.v(605)
    wire wand_781;   // mult.v(606)
    wire wand_812;   // mult.v(607)
    wire wand_843;   // mult.v(608)
    wire wfa_s_138;   // mult.v(609)
    wire wfa_cout_138;   // mult.v(609)
    wire wand_874;   // mult.v(610)
    wire wand_905;   // mult.v(611)
    wire wand_936;   // mult.v(612)
    wire wfa_s_139;   // mult.v(613)
    wire wfa_cout_139;   // mult.v(613)
    wire wand_255;   // mult.v(614)
    wire wand_286;   // mult.v(615)
    wire wand_317;   // mult.v(616)
    wire wfa_s_140;   // mult.v(617)
    wire wfa_cout_140;   // mult.v(617)
    wire wand_348;   // mult.v(618)
    wire wand_379;   // mult.v(619)
    wire wand_410;   // mult.v(620)
    wire wfa_s_141;   // mult.v(621)
    wire wfa_cout_141;   // mult.v(621)
    wire wand_441;   // mult.v(622)
    wire wand_472;   // mult.v(623)
    wire wand_503;   // mult.v(624)
    wire wfa_s_142;   // mult.v(625)
    wire wfa_cout_142;   // mult.v(625)
    wire wand_534;   // mult.v(626)
    wire wand_565;   // mult.v(627)
    wire wand_596;   // mult.v(628)
    wire wfa_s_143;   // mult.v(629)
    wire wfa_cout_143;   // mult.v(629)
    wire wand_627;   // mult.v(630)
    wire wand_658;   // mult.v(631)
    wire wand_689;   // mult.v(632)
    wire wfa_s_144;   // mult.v(633)
    wire wfa_cout_144;   // mult.v(633)
    wire wand_720;   // mult.v(634)
    wire wand_751;   // mult.v(635)
    wire wand_782;   // mult.v(636)
    wire wfa_s_145;   // mult.v(637)
    wire wfa_cout_145;   // mult.v(637)
    wire wand_813;   // mult.v(638)
    wire wand_844;   // mult.v(639)
    wire wand_875;   // mult.v(640)
    wire wfa_s_146;   // mult.v(641)
    wire wfa_cout_146;   // mult.v(641)
    wire wand_287;   // mult.v(642)
    wire wand_318;   // mult.v(643)
    wire wand_349;   // mult.v(644)
    wire wfa_s_147;   // mult.v(645)
    wire wfa_cout_147;   // mult.v(645)
    wire wand_380;   // mult.v(646)
    wire wand_411;   // mult.v(647)
    wire wand_442;   // mult.v(648)
    wire wfa_s_148;   // mult.v(649)
    wire wfa_cout_148;   // mult.v(649)
    wire wand_473;   // mult.v(650)
    wire wand_504;   // mult.v(651)
    wire wand_535;   // mult.v(652)
    wire wfa_s_149;   // mult.v(653)
    wire wfa_cout_149;   // mult.v(653)
    wire wand_566;   // mult.v(654)
    wire wand_597;   // mult.v(655)
    wire wand_628;   // mult.v(656)
    wire wfa_s_150;   // mult.v(657)
    wire wfa_cout_150;   // mult.v(657)
    wire wand_659;   // mult.v(658)
    wire wand_690;   // mult.v(659)
    wire wand_721;   // mult.v(660)
    wire wfa_s_151;   // mult.v(661)
    wire wfa_cout_151;   // mult.v(661)
    wire wand_752;   // mult.v(662)
    wire wand_783;   // mult.v(663)
    wire wand_814;   // mult.v(664)
    wire wfa_s_152;   // mult.v(665)
    wire wfa_cout_152;   // mult.v(665)
    wire wand_319;   // mult.v(666)
    wire wand_350;   // mult.v(667)
    wire wand_381;   // mult.v(668)
    wire wfa_s_153;   // mult.v(669)
    wire wfa_cout_153;   // mult.v(669)
    wire wand_412;   // mult.v(670)
    wire wand_443;   // mult.v(671)
    wire wand_474;   // mult.v(672)
    wire wfa_s_154;   // mult.v(673)
    wire wfa_cout_154;   // mult.v(673)
    wire wand_505;   // mult.v(674)
    wire wand_536;   // mult.v(675)
    wire wand_567;   // mult.v(676)
    wire wfa_s_155;   // mult.v(677)
    wire wfa_cout_155;   // mult.v(677)
    wire wand_598;   // mult.v(678)
    wire wand_629;   // mult.v(679)
    wire wand_660;   // mult.v(680)
    wire wfa_s_156;   // mult.v(681)
    wire wfa_cout_156;   // mult.v(681)
    wire wand_691;   // mult.v(682)
    wire wand_722;   // mult.v(683)
    wire wand_753;   // mult.v(684)
    wire wfa_s_157;   // mult.v(685)
    wire wfa_cout_157;   // mult.v(685)
    wire wand_351;   // mult.v(686)
    wire wand_382;   // mult.v(687)
    wire wand_413;   // mult.v(688)
    wire wfa_s_158;   // mult.v(689)
    wire wfa_cout_158;   // mult.v(689)
    wire wand_444;   // mult.v(690)
    wire wand_475;   // mult.v(691)
    wire wand_506;   // mult.v(692)
    wire wfa_s_159;   // mult.v(693)
    wire wfa_cout_159;   // mult.v(693)
    wire wand_537;   // mult.v(694)
    wire wand_568;   // mult.v(695)
    wire wand_599;   // mult.v(696)
    wire wfa_s_160;   // mult.v(697)
    wire wfa_cout_160;   // mult.v(697)
    wire wand_630;   // mult.v(698)
    wire wand_661;   // mult.v(699)
    wire wand_692;   // mult.v(700)
    wire wfa_s_161;   // mult.v(701)
    wire wfa_cout_161;   // mult.v(701)
    wire wand_383;   // mult.v(702)
    wire wand_414;   // mult.v(703)
    wire wand_445;   // mult.v(704)
    wire wfa_s_162;   // mult.v(705)
    wire wfa_cout_162;   // mult.v(705)
    wire wand_476;   // mult.v(706)
    wire wand_507;   // mult.v(707)
    wire wand_538;   // mult.v(708)
    wire wfa_s_163;   // mult.v(709)
    wire wfa_cout_163;   // mult.v(709)
    wire wand_569;   // mult.v(710)
    wire wand_600;   // mult.v(711)
    wire wand_631;   // mult.v(712)
    wire wfa_s_164;   // mult.v(713)
    wire wfa_cout_164;   // mult.v(713)
    wire wand_415;   // mult.v(714)
    wire wand_446;   // mult.v(715)
    wire wand_477;   // mult.v(716)
    wire wfa_s_165;   // mult.v(717)
    wire wfa_cout_165;   // mult.v(717)
    wire wand_508;   // mult.v(718)
    wire wand_539;   // mult.v(719)
    wire wand_570;   // mult.v(720)
    wire wfa_s_166;   // mult.v(721)
    wire wfa_cout_166;   // mult.v(721)
    wire wand_447;   // mult.v(722)
    wire wand_478;   // mult.v(723)
    wire wand_509;   // mult.v(724)
    wire wfa_s_167;   // mult.v(725)
    wire wfa_cout_167;   // mult.v(725)
    wire wand_13;   // mult.v(726)
    wire wand_44;   // mult.v(727)
    wire wha_s_14;   // mult.v(728)
    wire wha_c_14;   // mult.v(728)
    wire wand_14;   // mult.v(729)
    wire wand_45;   // mult.v(730)
    wire wand_76;   // mult.v(731)
    wire wfa_s_168;   // mult.v(732)
    wire wfa_cout_168;   // mult.v(732)
    wire wand_107;   // mult.v(733)
    wire wand_138;   // mult.v(734)
    wire wha_s_15;   // mult.v(735)
    wire wha_c_15;   // mult.v(735)
    wire wand_15;   // mult.v(736)
    wire wand_46;   // mult.v(737)
    wire wand_77;   // mult.v(738)
    wire wfa_s_169;   // mult.v(739)
    wire wfa_cout_169;   // mult.v(739)
    wire wand_108;   // mult.v(740)
    wire wand_139;   // mult.v(741)
    wire wand_170;   // mult.v(742)
    wire wfa_s_170;   // mult.v(743)
    wire wfa_cout_170;   // mult.v(743)
    wire wand_201;   // mult.v(744)
    wire wand_232;   // mult.v(745)
    wire wha_s_16;   // mult.v(746)
    wire wha_c_16;   // mult.v(746)
    wire wand_16;   // mult.v(747)
    wire wand_47;   // mult.v(748)
    wire wand_78;   // mult.v(749)
    wire wfa_s_171;   // mult.v(750)
    wire wfa_cout_171;   // mult.v(750)
    wire wand_109;   // mult.v(751)
    wire wand_140;   // mult.v(752)
    wire wand_171;   // mult.v(753)
    wire wfa_s_172;   // mult.v(754)
    wire wfa_cout_172;   // mult.v(754)
    wire wand_202;   // mult.v(755)
    wire wand_233;   // mult.v(756)
    wire wand_264;   // mult.v(757)
    wire wfa_s_173;   // mult.v(758)
    wire wfa_cout_173;   // mult.v(758)
    wire wand_295;   // mult.v(759)
    wire wand_326;   // mult.v(760)
    wire wha_s_17;   // mult.v(761)
    wire wha_c_17;   // mult.v(761)
    wire wand_17;   // mult.v(762)
    wire wand_48;   // mult.v(763)
    wire wand_79;   // mult.v(764)
    wire wfa_s_174;   // mult.v(765)
    wire wfa_cout_174;   // mult.v(765)
    wire wand_110;   // mult.v(766)
    wire wand_141;   // mult.v(767)
    wire wand_172;   // mult.v(768)
    wire wfa_s_175;   // mult.v(769)
    wire wfa_cout_175;   // mult.v(769)
    wire wand_203;   // mult.v(770)
    wire wand_234;   // mult.v(771)
    wire wand_265;   // mult.v(772)
    wire wfa_s_176;   // mult.v(773)
    wire wfa_cout_176;   // mult.v(773)
    wire wand_296;   // mult.v(774)
    wire wand_327;   // mult.v(775)
    wire wand_358;   // mult.v(776)
    wire wfa_s_177;   // mult.v(777)
    wire wfa_cout_177;   // mult.v(777)
    wire wand_389;   // mult.v(778)
    wire wand_420;   // mult.v(779)
    wire wha_s_18;   // mult.v(780)
    wire wha_c_18;   // mult.v(780)
    wire wand_18;   // mult.v(781)
    wire wand_49;   // mult.v(782)
    wire wand_80;   // mult.v(783)
    wire wfa_s_178;   // mult.v(784)
    wire wfa_cout_178;   // mult.v(784)
    wire wand_111;   // mult.v(785)
    wire wand_142;   // mult.v(786)
    wire wand_173;   // mult.v(787)
    wire wfa_s_179;   // mult.v(788)
    wire wfa_cout_179;   // mult.v(788)
    wire wand_204;   // mult.v(789)
    wire wand_235;   // mult.v(790)
    wire wand_266;   // mult.v(791)
    wire wfa_s_180;   // mult.v(792)
    wire wfa_cout_180;   // mult.v(792)
    wire wand_297;   // mult.v(793)
    wire wand_328;   // mult.v(794)
    wire wand_359;   // mult.v(795)
    wire wfa_s_181;   // mult.v(796)
    wire wfa_cout_181;   // mult.v(796)
    wire wand_390;   // mult.v(797)
    wire wand_421;   // mult.v(798)
    wire wand_452;   // mult.v(799)
    wire wfa_s_182;   // mult.v(800)
    wire wfa_cout_182;   // mult.v(800)
    wire wand_483;   // mult.v(801)
    wire wand_514;   // mult.v(802)
    wire wha_s_19;   // mult.v(803)
    wire wha_c_19;   // mult.v(803)
    wire wand_81;   // mult.v(804)
    wire wand_112;   // mult.v(805)
    wire wand_143;   // mult.v(806)
    wire wfa_s_183;   // mult.v(807)
    wire wfa_cout_183;   // mult.v(807)
    wire wand_174;   // mult.v(808)
    wire wand_205;   // mult.v(809)
    wire wand_236;   // mult.v(810)
    wire wfa_s_184;   // mult.v(811)
    wire wfa_cout_184;   // mult.v(811)
    wire wand_267;   // mult.v(812)
    wire wand_298;   // mult.v(813)
    wire wand_329;   // mult.v(814)
    wire wfa_s_185;   // mult.v(815)
    wire wfa_cout_185;   // mult.v(815)
    wire wand_360;   // mult.v(816)
    wire wand_391;   // mult.v(817)
    wire wand_422;   // mult.v(818)
    wire wfa_s_186;   // mult.v(819)
    wire wfa_cout_186;   // mult.v(819)
    wire wand_453;   // mult.v(820)
    wire wand_484;   // mult.v(821)
    wire wand_515;   // mult.v(822)
    wire wfa_s_187;   // mult.v(823)
    wire wfa_cout_187;   // mult.v(823)
    wire wand_546;   // mult.v(824)
    wire wand_577;   // mult.v(825)
    wire wand_608;   // mult.v(826)
    wire wfa_s_188;   // mult.v(827)
    wire wfa_cout_188;   // mult.v(827)
    wire wand_175;   // mult.v(828)
    wire wand_206;   // mult.v(829)
    wire wand_237;   // mult.v(830)
    wire wfa_s_189;   // mult.v(831)
    wire wfa_cout_189;   // mult.v(831)
    wire wand_268;   // mult.v(832)
    wire wand_299;   // mult.v(833)
    wire wand_330;   // mult.v(834)
    wire wfa_s_190;   // mult.v(835)
    wire wfa_cout_190;   // mult.v(835)
    wire wand_361;   // mult.v(836)
    wire wand_392;   // mult.v(837)
    wire wand_423;   // mult.v(838)
    wire wfa_s_191;   // mult.v(839)
    wire wfa_cout_191;   // mult.v(839)
    wire wand_454;   // mult.v(840)
    wire wand_485;   // mult.v(841)
    wire wand_516;   // mult.v(842)
    wire wfa_s_192;   // mult.v(843)
    wire wfa_cout_192;   // mult.v(843)
    wire wand_547;   // mult.v(844)
    wire wand_578;   // mult.v(845)
    wire wand_609;   // mult.v(846)
    wire wfa_s_193;   // mult.v(847)
    wire wfa_cout_193;   // mult.v(847)
    wire wand_640;   // mult.v(848)
    wire wfa_s_194;   // mult.v(849)
    wire wfa_cout_194;   // mult.v(849)
    wire wand_269;   // mult.v(850)
    wire wand_300;   // mult.v(851)
    wire wand_331;   // mult.v(852)
    wire wfa_s_195;   // mult.v(853)
    wire wfa_cout_195;   // mult.v(853)
    wire wand_362;   // mult.v(854)
    wire wand_393;   // mult.v(855)
    wire wand_424;   // mult.v(856)
    wire wfa_s_196;   // mult.v(857)
    wire wfa_cout_196;   // mult.v(857)
    wire wand_455;   // mult.v(858)
    wire wand_486;   // mult.v(859)
    wire wand_517;   // mult.v(860)
    wire wfa_s_197;   // mult.v(861)
    wire wfa_cout_197;   // mult.v(861)
    wire wand_548;   // mult.v(862)
    wire wand_579;   // mult.v(863)
    wire wand_610;   // mult.v(864)
    wire wfa_s_198;   // mult.v(865)
    wire wfa_cout_198;   // mult.v(865)
    wire wand_641;   // mult.v(866)
    wire wand_672;   // mult.v(867)
    wire wfa_s_199;   // mult.v(868)
    wire wfa_cout_199;   // mult.v(868)
    wire wfa_s_200;   // mult.v(869)
    wire wfa_cout_200;   // mult.v(869)
    wire wand_363;   // mult.v(870)
    wire wand_394;   // mult.v(871)
    wire wand_425;   // mult.v(872)
    wire wfa_s_201;   // mult.v(873)
    wire wfa_cout_201;   // mult.v(873)
    wire wand_456;   // mult.v(874)
    wire wand_487;   // mult.v(875)
    wire wand_518;   // mult.v(876)
    wire wfa_s_202;   // mult.v(877)
    wire wfa_cout_202;   // mult.v(877)
    wire wand_549;   // mult.v(878)
    wire wand_580;   // mult.v(879)
    wire wand_611;   // mult.v(880)
    wire wfa_s_203;   // mult.v(881)
    wire wfa_cout_203;   // mult.v(881)
    wire wand_642;   // mult.v(882)
    wire wand_673;   // mult.v(883)
    wire wand_704;   // mult.v(884)
    wire wfa_s_204;   // mult.v(885)
    wire wfa_cout_204;   // mult.v(885)
    wire wfa_s_205;   // mult.v(886)
    wire wfa_cout_205;   // mult.v(886)
    wire wfa_s_206;   // mult.v(887)
    wire wfa_cout_206;   // mult.v(887)
    wire wand_457;   // mult.v(888)
    wire wand_488;   // mult.v(889)
    wire wand_519;   // mult.v(890)
    wire wfa_s_207;   // mult.v(891)
    wire wfa_cout_207;   // mult.v(891)
    wire wand_550;   // mult.v(892)
    wire wand_581;   // mult.v(893)
    wire wand_612;   // mult.v(894)
    wire wfa_s_208;   // mult.v(895)
    wire wfa_cout_208;   // mult.v(895)
    wire wand_643;   // mult.v(896)
    wire wand_674;   // mult.v(897)
    wire wand_705;   // mult.v(898)
    wire wfa_s_209;   // mult.v(899)
    wire wfa_cout_209;   // mult.v(899)
    wire wand_736;   // mult.v(900)
    wire wfa_s_210;   // mult.v(901)
    wire wfa_cout_210;   // mult.v(901)
    wire wfa_s_211;   // mult.v(902)
    wire wfa_cout_211;   // mult.v(902)
    wire wfa_s_212;   // mult.v(903)
    wire wfa_cout_212;   // mult.v(903)
    wire wand_551;   // mult.v(904)
    wire wand_582;   // mult.v(905)
    wire wand_613;   // mult.v(906)
    wire wfa_s_213;   // mult.v(907)
    wire wfa_cout_213;   // mult.v(907)
    wire wand_644;   // mult.v(908)
    wire wand_675;   // mult.v(909)
    wire wand_706;   // mult.v(910)
    wire wfa_s_214;   // mult.v(911)
    wire wfa_cout_214;   // mult.v(911)
    wire wand_737;   // mult.v(912)
    wire wand_768;   // mult.v(913)
    wire wfa_s_215;   // mult.v(914)
    wire wfa_cout_215;   // mult.v(914)
    wire wfa_s_216;   // mult.v(915)
    wire wfa_cout_216;   // mult.v(915)
    wire wfa_s_217;   // mult.v(916)
    wire wfa_cout_217;   // mult.v(916)
    wire wfa_s_218;   // mult.v(917)
    wire wfa_cout_218;   // mult.v(917)
    wire wand_645;   // mult.v(918)
    wire wand_676;   // mult.v(919)
    wire wand_707;   // mult.v(920)
    wire wfa_s_219;   // mult.v(921)
    wire wfa_cout_219;   // mult.v(921)
    wire wand_738;   // mult.v(922)
    wire wand_769;   // mult.v(923)
    wire wand_800;   // mult.v(924)
    wire wfa_s_220;   // mult.v(925)
    wire wfa_cout_220;   // mult.v(925)
    wire wfa_s_221;   // mult.v(926)
    wire wfa_cout_221;   // mult.v(926)
    wire wfa_s_222;   // mult.v(927)
    wire wfa_cout_222;   // mult.v(927)
    wire wfa_s_223;   // mult.v(928)
    wire wfa_cout_223;   // mult.v(928)
    wire wfa_s_224;   // mult.v(929)
    wire wfa_cout_224;   // mult.v(929)
    wire wand_739;   // mult.v(930)
    wire wand_770;   // mult.v(931)
    wire wand_801;   // mult.v(932)
    wire wfa_s_225;   // mult.v(933)
    wire wfa_cout_225;   // mult.v(933)
    wire wand_832;   // mult.v(934)
    wire wfa_s_226;   // mult.v(935)
    wire wfa_cout_226;   // mult.v(935)
    wire wfa_s_227;   // mult.v(936)
    wire wfa_cout_227;   // mult.v(936)
    wire wfa_s_228;   // mult.v(937)
    wire wfa_cout_228;   // mult.v(937)
    wire wfa_s_229;   // mult.v(938)
    wire wfa_cout_229;   // mult.v(938)
    wire wfa_s_230;   // mult.v(939)
    wire wfa_cout_230;   // mult.v(939)
    wire wand_833;   // mult.v(940)
    wire wand_864;   // mult.v(941)
    wire wfa_s_231;   // mult.v(942)
    wire wfa_cout_231;   // mult.v(942)
    wire wfa_s_232;   // mult.v(943)
    wire wfa_cout_232;   // mult.v(943)
    wire wfa_s_233;   // mult.v(944)
    wire wfa_cout_233;   // mult.v(944)
    wire wfa_s_234;   // mult.v(945)
    wire wfa_cout_234;   // mult.v(945)
    wire wfa_s_235;   // mult.v(946)
    wire wfa_cout_235;   // mult.v(946)
    wire wfa_s_236;   // mult.v(947)
    wire wfa_cout_236;   // mult.v(947)
    wire wfa_s_237;   // mult.v(948)
    wire wfa_cout_237;   // mult.v(948)
    wire wfa_s_238;   // mult.v(949)
    wire wfa_cout_238;   // mult.v(949)
    wire wfa_s_239;   // mult.v(950)
    wire wfa_cout_239;   // mult.v(950)
    wire wfa_s_240;   // mult.v(951)
    wire wfa_cout_240;   // mult.v(951)
    wire wfa_s_241;   // mult.v(952)
    wire wfa_cout_241;   // mult.v(952)
    wire wfa_s_242;   // mult.v(953)
    wire wfa_cout_242;   // mult.v(953)
    wire wfa_s_243;   // mult.v(954)
    wire wfa_cout_243;   // mult.v(954)
    wire wfa_s_244;   // mult.v(955)
    wire wfa_cout_244;   // mult.v(955)
    wire wfa_s_245;   // mult.v(956)
    wire wfa_cout_245;   // mult.v(956)
    wire wfa_s_246;   // mult.v(957)
    wire wfa_cout_246;   // mult.v(957)
    wire wfa_s_247;   // mult.v(958)
    wire wfa_cout_247;   // mult.v(958)
    wire wfa_s_248;   // mult.v(959)
    wire wfa_cout_248;   // mult.v(959)
    wire wfa_s_249;   // mult.v(960)
    wire wfa_cout_249;   // mult.v(960)
    wire wfa_s_250;   // mult.v(961)
    wire wfa_cout_250;   // mult.v(961)
    wire wfa_s_251;   // mult.v(962)
    wire wfa_cout_251;   // mult.v(962)
    wire wfa_s_252;   // mult.v(963)
    wire wfa_cout_252;   // mult.v(963)
    wire wfa_s_253;   // mult.v(964)
    wire wfa_cout_253;   // mult.v(964)
    wire wfa_s_254;   // mult.v(965)
    wire wfa_cout_254;   // mult.v(965)
    wire wfa_s_255;   // mult.v(966)
    wire wfa_cout_255;   // mult.v(966)
    wire wfa_s_256;   // mult.v(967)
    wire wfa_cout_256;   // mult.v(967)
    wire wfa_s_257;   // mult.v(968)
    wire wfa_cout_257;   // mult.v(968)
    wire wfa_s_258;   // mult.v(969)
    wire wfa_cout_258;   // mult.v(969)
    wire wfa_s_259;   // mult.v(970)
    wire wfa_cout_259;   // mult.v(970)
    wire wfa_s_260;   // mult.v(971)
    wire wfa_cout_260;   // mult.v(971)
    wire wfa_s_261;   // mult.v(972)
    wire wfa_cout_261;   // mult.v(972)
    wire wfa_s_262;   // mult.v(973)
    wire wfa_cout_262;   // mult.v(973)
    wire wfa_s_263;   // mult.v(974)
    wire wfa_cout_263;   // mult.v(974)
    wire wfa_s_264;   // mult.v(975)
    wire wfa_cout_264;   // mult.v(975)
    wire wfa_s_265;   // mult.v(976)
    wire wfa_cout_265;   // mult.v(976)
    wire wfa_s_266;   // mult.v(977)
    wire wfa_cout_266;   // mult.v(977)
    wire wfa_s_267;   // mult.v(978)
    wire wfa_cout_267;   // mult.v(978)
    wire wfa_s_268;   // mult.v(979)
    wire wfa_cout_268;   // mult.v(979)
    wire wfa_s_269;   // mult.v(980)
    wire wfa_cout_269;   // mult.v(980)
    wire wfa_s_270;   // mult.v(981)
    wire wfa_cout_270;   // mult.v(981)
    wire wfa_s_271;   // mult.v(982)
    wire wfa_cout_271;   // mult.v(982)
    wire wfa_s_272;   // mult.v(983)
    wire wfa_cout_272;   // mult.v(983)
    wire wfa_s_273;   // mult.v(984)
    wire wfa_cout_273;   // mult.v(984)
    wire wfa_s_274;   // mult.v(985)
    wire wfa_cout_274;   // mult.v(985)
    wire wfa_s_275;   // mult.v(986)
    wire wfa_cout_275;   // mult.v(986)
    wire wfa_s_276;   // mult.v(987)
    wire wfa_cout_276;   // mult.v(987)
    wire wfa_s_277;   // mult.v(988)
    wire wfa_cout_277;   // mult.v(988)
    wire wfa_s_278;   // mult.v(989)
    wire wfa_cout_278;   // mult.v(989)
    wire wfa_s_279;   // mult.v(990)
    wire wfa_cout_279;   // mult.v(990)
    wire wfa_s_280;   // mult.v(991)
    wire wfa_cout_280;   // mult.v(991)
    wire wfa_s_281;   // mult.v(992)
    wire wfa_cout_281;   // mult.v(992)
    wire wfa_s_282;   // mult.v(993)
    wire wfa_cout_282;   // mult.v(993)
    wire wfa_s_283;   // mult.v(994)
    wire wfa_cout_283;   // mult.v(994)
    wire wfa_s_284;   // mult.v(995)
    wire wfa_cout_284;   // mult.v(995)
    wire wfa_s_285;   // mult.v(996)
    wire wfa_cout_285;   // mult.v(996)
    wire wfa_s_286;   // mult.v(997)
    wire wfa_cout_286;   // mult.v(997)
    wire wfa_s_287;   // mult.v(998)
    wire wfa_cout_287;   // mult.v(998)
    wire wfa_s_288;   // mult.v(999)
    wire wfa_cout_288;   // mult.v(999)
    wire wfa_s_289;   // mult.v(1000)
    wire wfa_cout_289;   // mult.v(1000)
    wire wfa_s_290;   // mult.v(1001)
    wire wfa_cout_290;   // mult.v(1001)
    wire wand_967;   // mult.v(1002)
    wire wand_998;   // mult.v(1003)
    wire wfa_s_291;   // mult.v(1004)
    wire wfa_cout_291;   // mult.v(1004)
    wire wfa_s_292;   // mult.v(1005)
    wire wfa_cout_292;   // mult.v(1005)
    wire wfa_s_293;   // mult.v(1006)
    wire wfa_cout_293;   // mult.v(1006)
    wire wfa_s_294;   // mult.v(1007)
    wire wfa_cout_294;   // mult.v(1007)
    wire wfa_s_295;   // mult.v(1008)
    wire wfa_cout_295;   // mult.v(1008)
    wire wfa_s_296;   // mult.v(1009)
    wire wfa_cout_296;   // mult.v(1009)
    wire wand_906;   // mult.v(1010)
    wire wand_937;   // mult.v(1011)
    wire wand_968;   // mult.v(1012)
    wire wfa_s_297;   // mult.v(1013)
    wire wfa_cout_297;   // mult.v(1013)
    wire wand_999;   // mult.v(1014)
    wire wfa_s_298;   // mult.v(1015)
    wire wfa_cout_298;   // mult.v(1015)
    wire wfa_s_299;   // mult.v(1016)
    wire wfa_cout_299;   // mult.v(1016)
    wire wfa_s_300;   // mult.v(1017)
    wire wfa_cout_300;   // mult.v(1017)
    wire wfa_s_301;   // mult.v(1018)
    wire wfa_cout_301;   // mult.v(1018)
    wire wfa_s_302;   // mult.v(1019)
    wire wfa_cout_302;   // mult.v(1019)
    wire wand_845;   // mult.v(1020)
    wire wand_876;   // mult.v(1021)
    wire wand_907;   // mult.v(1022)
    wire wfa_s_303;   // mult.v(1023)
    wire wfa_cout_303;   // mult.v(1023)
    wire wand_938;   // mult.v(1024)
    wire wand_969;   // mult.v(1025)
    wire wand_1000;   // mult.v(1026)
    wire wfa_s_304;   // mult.v(1027)
    wire wfa_cout_304;   // mult.v(1027)
    wire wfa_s_305;   // mult.v(1028)
    wire wfa_cout_305;   // mult.v(1028)
    wire wfa_s_306;   // mult.v(1029)
    wire wfa_cout_306;   // mult.v(1029)
    wire wfa_s_307;   // mult.v(1030)
    wire wfa_cout_307;   // mult.v(1030)
    wire wfa_s_308;   // mult.v(1031)
    wire wfa_cout_308;   // mult.v(1031)
    wire wand_784;   // mult.v(1032)
    wire wand_815;   // mult.v(1033)
    wire wand_846;   // mult.v(1034)
    wire wfa_s_309;   // mult.v(1035)
    wire wfa_cout_309;   // mult.v(1035)
    wire wand_877;   // mult.v(1036)
    wire wand_908;   // mult.v(1037)
    wire wand_939;   // mult.v(1038)
    wire wfa_s_310;   // mult.v(1039)
    wire wfa_cout_310;   // mult.v(1039)
    wire wand_970;   // mult.v(1040)
    wire wand_1001;   // mult.v(1041)
    wire wfa_s_311;   // mult.v(1042)
    wire wfa_cout_311;   // mult.v(1042)
    wire wfa_s_312;   // mult.v(1043)
    wire wfa_cout_312;   // mult.v(1043)
    wire wfa_s_313;   // mult.v(1044)
    wire wfa_cout_313;   // mult.v(1044)
    wire wfa_s_314;   // mult.v(1045)
    wire wfa_cout_314;   // mult.v(1045)
    wire wand_723;   // mult.v(1046)
    wire wand_754;   // mult.v(1047)
    wire wand_785;   // mult.v(1048)
    wire wfa_s_315;   // mult.v(1049)
    wire wfa_cout_315;   // mult.v(1049)
    wire wand_816;   // mult.v(1050)
    wire wand_847;   // mult.v(1051)
    wire wand_878;   // mult.v(1052)
    wire wfa_s_316;   // mult.v(1053)
    wire wfa_cout_316;   // mult.v(1053)
    wire wand_909;   // mult.v(1054)
    wire wand_940;   // mult.v(1055)
    wire wand_971;   // mult.v(1056)
    wire wfa_s_317;   // mult.v(1057)
    wire wfa_cout_317;   // mult.v(1057)
    wire wand_1002;   // mult.v(1058)
    wire wfa_s_318;   // mult.v(1059)
    wire wfa_cout_318;   // mult.v(1059)
    wire wfa_s_319;   // mult.v(1060)
    wire wfa_cout_319;   // mult.v(1060)
    wire wfa_s_320;   // mult.v(1061)
    wire wfa_cout_320;   // mult.v(1061)
    wire wand_662;   // mult.v(1062)
    wire wand_693;   // mult.v(1063)
    wire wand_724;   // mult.v(1064)
    wire wfa_s_321;   // mult.v(1065)
    wire wfa_cout_321;   // mult.v(1065)
    wire wand_755;   // mult.v(1066)
    wire wand_786;   // mult.v(1067)
    wire wand_817;   // mult.v(1068)
    wire wfa_s_322;   // mult.v(1069)
    wire wfa_cout_322;   // mult.v(1069)
    wire wand_848;   // mult.v(1070)
    wire wand_879;   // mult.v(1071)
    wire wand_910;   // mult.v(1072)
    wire wfa_s_323;   // mult.v(1073)
    wire wfa_cout_323;   // mult.v(1073)
    wire wand_941;   // mult.v(1074)
    wire wand_972;   // mult.v(1075)
    wire wand_1003;   // mult.v(1076)
    wire wfa_s_324;   // mult.v(1077)
    wire wfa_cout_324;   // mult.v(1077)
    wire wfa_s_325;   // mult.v(1078)
    wire wfa_cout_325;   // mult.v(1078)
    wire wfa_s_326;   // mult.v(1079)
    wire wfa_cout_326;   // mult.v(1079)
    wire wand_601;   // mult.v(1080)
    wire wand_632;   // mult.v(1081)
    wire wand_663;   // mult.v(1082)
    wire wfa_s_327;   // mult.v(1083)
    wire wfa_cout_327;   // mult.v(1083)
    wire wand_694;   // mult.v(1084)
    wire wand_725;   // mult.v(1085)
    wire wand_756;   // mult.v(1086)
    wire wfa_s_328;   // mult.v(1087)
    wire wfa_cout_328;   // mult.v(1087)
    wire wand_787;   // mult.v(1088)
    wire wand_818;   // mult.v(1089)
    wire wand_849;   // mult.v(1090)
    wire wfa_s_329;   // mult.v(1091)
    wire wfa_cout_329;   // mult.v(1091)
    wire wand_880;   // mult.v(1092)
    wire wand_911;   // mult.v(1093)
    wire wand_942;   // mult.v(1094)
    wire wfa_s_330;   // mult.v(1095)
    wire wfa_cout_330;   // mult.v(1095)
    wire wand_973;   // mult.v(1096)
    wire wand_1004;   // mult.v(1097)
    wire wfa_s_331;   // mult.v(1098)
    wire wfa_cout_331;   // mult.v(1098)
    wire wfa_s_332;   // mult.v(1099)
    wire wfa_cout_332;   // mult.v(1099)
    wire wand_540;   // mult.v(1100)
    wire wand_571;   // mult.v(1101)
    wire wand_602;   // mult.v(1102)
    wire wfa_s_333;   // mult.v(1103)
    wire wfa_cout_333;   // mult.v(1103)
    wire wand_633;   // mult.v(1104)
    wire wand_664;   // mult.v(1105)
    wire wand_695;   // mult.v(1106)
    wire wfa_s_334;   // mult.v(1107)
    wire wfa_cout_334;   // mult.v(1107)
    wire wand_726;   // mult.v(1108)
    wire wand_757;   // mult.v(1109)
    wire wand_788;   // mult.v(1110)
    wire wfa_s_335;   // mult.v(1111)
    wire wfa_cout_335;   // mult.v(1111)
    wire wand_819;   // mult.v(1112)
    wire wand_850;   // mult.v(1113)
    wire wand_881;   // mult.v(1114)
    wire wfa_s_336;   // mult.v(1115)
    wire wfa_cout_336;   // mult.v(1115)
    wire wand_912;   // mult.v(1116)
    wire wand_943;   // mult.v(1117)
    wire wand_974;   // mult.v(1118)
    wire wfa_s_337;   // mult.v(1119)
    wire wfa_cout_337;   // mult.v(1119)
    wire wand_1005;   // mult.v(1120)
    wire wfa_s_338;   // mult.v(1121)
    wire wfa_cout_338;   // mult.v(1121)
    wire wand_479;   // mult.v(1122)
    wire wand_510;   // mult.v(1123)
    wire wand_541;   // mult.v(1124)
    wire wfa_s_339;   // mult.v(1125)
    wire wfa_cout_339;   // mult.v(1125)
    wire wand_572;   // mult.v(1126)
    wire wand_603;   // mult.v(1127)
    wire wand_634;   // mult.v(1128)
    wire wfa_s_340;   // mult.v(1129)
    wire wfa_cout_340;   // mult.v(1129)
    wire wand_665;   // mult.v(1130)
    wire wand_696;   // mult.v(1131)
    wire wand_727;   // mult.v(1132)
    wire wfa_s_341;   // mult.v(1133)
    wire wfa_cout_341;   // mult.v(1133)
    wire wand_758;   // mult.v(1134)
    wire wand_789;   // mult.v(1135)
    wire wand_820;   // mult.v(1136)
    wire wfa_s_342;   // mult.v(1137)
    wire wfa_cout_342;   // mult.v(1137)
    wire wand_851;   // mult.v(1138)
    wire wand_882;   // mult.v(1139)
    wire wand_913;   // mult.v(1140)
    wire wfa_s_343;   // mult.v(1141)
    wire wfa_cout_343;   // mult.v(1141)
    wire wand_944;   // mult.v(1142)
    wire wand_975;   // mult.v(1143)
    wire wand_1006;   // mult.v(1144)
    wire wfa_s_344;   // mult.v(1145)
    wire wfa_cout_344;   // mult.v(1145)
    wire wand_511;   // mult.v(1146)
    wire wand_542;   // mult.v(1147)
    wire wand_573;   // mult.v(1148)
    wire wfa_s_345;   // mult.v(1149)
    wire wfa_cout_345;   // mult.v(1149)
    wire wand_604;   // mult.v(1150)
    wire wand_635;   // mult.v(1151)
    wire wand_666;   // mult.v(1152)
    wire wfa_s_346;   // mult.v(1153)
    wire wfa_cout_346;   // mult.v(1153)
    wire wand_697;   // mult.v(1154)
    wire wand_728;   // mult.v(1155)
    wire wand_759;   // mult.v(1156)
    wire wfa_s_347;   // mult.v(1157)
    wire wfa_cout_347;   // mult.v(1157)
    wire wand_790;   // mult.v(1158)
    wire wand_821;   // mult.v(1159)
    wire wand_852;   // mult.v(1160)
    wire wfa_s_348;   // mult.v(1161)
    wire wfa_cout_348;   // mult.v(1161)
    wire wand_883;   // mult.v(1162)
    wire wand_914;   // mult.v(1163)
    wire wand_945;   // mult.v(1164)
    wire wfa_s_349;   // mult.v(1165)
    wire wfa_cout_349;   // mult.v(1165)
    wire wand_543;   // mult.v(1166)
    wire wand_574;   // mult.v(1167)
    wire wand_605;   // mult.v(1168)
    wire wfa_s_350;   // mult.v(1169)
    wire wfa_cout_350;   // mult.v(1169)
    wire wand_636;   // mult.v(1170)
    wire wand_667;   // mult.v(1171)
    wire wand_698;   // mult.v(1172)
    wire wfa_s_351;   // mult.v(1173)
    wire wfa_cout_351;   // mult.v(1173)
    wire wand_729;   // mult.v(1174)
    wire wand_760;   // mult.v(1175)
    wire wand_791;   // mult.v(1176)
    wire wfa_s_352;   // mult.v(1177)
    wire wfa_cout_352;   // mult.v(1177)
    wire wand_822;   // mult.v(1178)
    wire wand_853;   // mult.v(1179)
    wire wand_884;   // mult.v(1180)
    wire wfa_s_353;   // mult.v(1181)
    wire wfa_cout_353;   // mult.v(1181)
    wire wand_575;   // mult.v(1182)
    wire wand_606;   // mult.v(1183)
    wire wand_637;   // mult.v(1184)
    wire wfa_s_354;   // mult.v(1185)
    wire wfa_cout_354;   // mult.v(1185)
    wire wand_668;   // mult.v(1186)
    wire wand_699;   // mult.v(1187)
    wire wand_730;   // mult.v(1188)
    wire wfa_s_355;   // mult.v(1189)
    wire wfa_cout_355;   // mult.v(1189)
    wire wand_761;   // mult.v(1190)
    wire wand_792;   // mult.v(1191)
    wire wand_823;   // mult.v(1192)
    wire wfa_s_356;   // mult.v(1193)
    wire wfa_cout_356;   // mult.v(1193)
    wire wand_607;   // mult.v(1194)
    wire wand_638;   // mult.v(1195)
    wire wand_669;   // mult.v(1196)
    wire wfa_s_357;   // mult.v(1197)
    wire wfa_cout_357;   // mult.v(1197)
    wire wand_700;   // mult.v(1198)
    wire wand_731;   // mult.v(1199)
    wire wand_762;   // mult.v(1200)
    wire wfa_s_358;   // mult.v(1201)
    wire wfa_cout_358;   // mult.v(1201)
    wire wand_639;   // mult.v(1202)
    wire wand_670;   // mult.v(1203)
    wire wand_701;   // mult.v(1204)
    wire wfa_s_359;   // mult.v(1205)
    wire wfa_cout_359;   // mult.v(1205)
    wire wand_9;   // mult.v(1206)
    wire wand_40;   // mult.v(1207)
    wire wha_s_20;   // mult.v(1208)
    wire wha_c_20;   // mult.v(1208)
    wire wand_10;   // mult.v(1209)
    wire wand_41;   // mult.v(1210)
    wire wand_72;   // mult.v(1211)
    wire wfa_s_360;   // mult.v(1212)
    wire wfa_cout_360;   // mult.v(1212)
    wire wand_103;   // mult.v(1213)
    wire wand_134;   // mult.v(1214)
    wire wha_s_21;   // mult.v(1215)
    wire wha_c_21;   // mult.v(1215)
    wire wand_11;   // mult.v(1216)
    wire wand_42;   // mult.v(1217)
    wire wand_73;   // mult.v(1218)
    wire wfa_s_361;   // mult.v(1219)
    wire wfa_cout_361;   // mult.v(1219)
    wire wand_104;   // mult.v(1220)
    wire wand_135;   // mult.v(1221)
    wire wand_166;   // mult.v(1222)
    wire wfa_s_362;   // mult.v(1223)
    wire wfa_cout_362;   // mult.v(1223)
    wire wand_197;   // mult.v(1224)
    wire wand_228;   // mult.v(1225)
    wire wha_s_22;   // mult.v(1226)
    wire wha_c_22;   // mult.v(1226)
    wire wand_12;   // mult.v(1227)
    wire wand_43;   // mult.v(1228)
    wire wand_74;   // mult.v(1229)
    wire wfa_s_363;   // mult.v(1230)
    wire wfa_cout_363;   // mult.v(1230)
    wire wand_105;   // mult.v(1231)
    wire wand_136;   // mult.v(1232)
    wire wand_167;   // mult.v(1233)
    wire wfa_s_364;   // mult.v(1234)
    wire wfa_cout_364;   // mult.v(1234)
    wire wand_198;   // mult.v(1235)
    wire wand_229;   // mult.v(1236)
    wire wand_260;   // mult.v(1237)
    wire wfa_s_365;   // mult.v(1238)
    wire wfa_cout_365;   // mult.v(1238)
    wire wand_291;   // mult.v(1239)
    wire wand_322;   // mult.v(1240)
    wire wha_s_23;   // mult.v(1241)
    wire wha_c_23;   // mult.v(1241)
    wire wand_75;   // mult.v(1242)
    wire wand_106;   // mult.v(1243)
    wire wand_137;   // mult.v(1244)
    wire wfa_s_366;   // mult.v(1245)
    wire wfa_cout_366;   // mult.v(1245)
    wire wand_168;   // mult.v(1246)
    wire wand_199;   // mult.v(1247)
    wire wand_230;   // mult.v(1248)
    wire wfa_s_367;   // mult.v(1249)
    wire wfa_cout_367;   // mult.v(1249)
    wire wand_261;   // mult.v(1250)
    wire wand_292;   // mult.v(1251)
    wire wand_323;   // mult.v(1252)
    wire wfa_s_368;   // mult.v(1253)
    wire wfa_cout_368;   // mult.v(1253)
    wire wand_354;   // mult.v(1254)
    wire wand_385;   // mult.v(1255)
    wire wand_416;   // mult.v(1256)
    wire wfa_s_369;   // mult.v(1257)
    wire wfa_cout_369;   // mult.v(1257)
    wire wand_169;   // mult.v(1258)
    wire wand_200;   // mult.v(1259)
    wire wand_231;   // mult.v(1260)
    wire wfa_s_370;   // mult.v(1261)
    wire wfa_cout_370;   // mult.v(1261)
    wire wand_262;   // mult.v(1262)
    wire wand_293;   // mult.v(1263)
    wire wand_324;   // mult.v(1264)
    wire wfa_s_371;   // mult.v(1265)
    wire wfa_cout_371;   // mult.v(1265)
    wire wand_355;   // mult.v(1266)
    wire wand_386;   // mult.v(1267)
    wire wand_417;   // mult.v(1268)
    wire wfa_s_372;   // mult.v(1269)
    wire wfa_cout_372;   // mult.v(1269)
    wire wand_448;   // mult.v(1270)
    wire wfa_s_373;   // mult.v(1271)
    wire wfa_cout_373;   // mult.v(1271)
    wire wand_263;   // mult.v(1272)
    wire wand_294;   // mult.v(1273)
    wire wand_325;   // mult.v(1274)
    wire wfa_s_374;   // mult.v(1275)
    wire wfa_cout_374;   // mult.v(1275)
    wire wand_356;   // mult.v(1276)
    wire wand_387;   // mult.v(1277)
    wire wand_418;   // mult.v(1278)
    wire wfa_s_375;   // mult.v(1279)
    wire wfa_cout_375;   // mult.v(1279)
    wire wand_449;   // mult.v(1280)
    wire wand_480;   // mult.v(1281)
    wire wfa_s_376;   // mult.v(1282)
    wire wfa_cout_376;   // mult.v(1282)
    wire wfa_s_377;   // mult.v(1283)
    wire wfa_cout_377;   // mult.v(1283)
    wire wand_357;   // mult.v(1284)
    wire wand_388;   // mult.v(1285)
    wire wand_419;   // mult.v(1286)
    wire wfa_s_378;   // mult.v(1287)
    wire wfa_cout_378;   // mult.v(1287)
    wire wand_450;   // mult.v(1288)
    wire wand_481;   // mult.v(1289)
    wire wand_512;   // mult.v(1290)
    wire wfa_s_379;   // mult.v(1291)
    wire wfa_cout_379;   // mult.v(1291)
    wire wfa_s_380;   // mult.v(1292)
    wire wfa_cout_380;   // mult.v(1292)
    wire wfa_s_381;   // mult.v(1293)
    wire wfa_cout_381;   // mult.v(1293)
    wire wand_451;   // mult.v(1294)
    wire wand_482;   // mult.v(1295)
    wire wand_513;   // mult.v(1296)
    wire wfa_s_382;   // mult.v(1297)
    wire wfa_cout_382;   // mult.v(1297)
    wire wand_544;   // mult.v(1298)
    wire wfa_s_383;   // mult.v(1299)
    wire wfa_cout_383;   // mult.v(1299)
    wire wfa_s_384;   // mult.v(1300)
    wire wfa_cout_384;   // mult.v(1300)
    wire wfa_s_385;   // mult.v(1301)
    wire wfa_cout_385;   // mult.v(1301)
    wire wand_545;   // mult.v(1302)
    wire wand_576;   // mult.v(1303)
    wire wfa_s_386;   // mult.v(1304)
    wire wfa_cout_386;   // mult.v(1304)
    wire wfa_s_387;   // mult.v(1305)
    wire wfa_cout_387;   // mult.v(1305)
    wire wfa_s_388;   // mult.v(1306)
    wire wfa_cout_388;   // mult.v(1306)
    wire wfa_s_389;   // mult.v(1307)
    wire wfa_cout_389;   // mult.v(1307)
    wire wfa_s_390;   // mult.v(1308)
    wire wfa_cout_390;   // mult.v(1308)
    wire wfa_s_391;   // mult.v(1309)
    wire wfa_cout_391;   // mult.v(1309)
    wire wfa_s_392;   // mult.v(1310)
    wire wfa_cout_392;   // mult.v(1310)
    wire wfa_s_393;   // mult.v(1311)
    wire wfa_cout_393;   // mult.v(1311)
    wire wfa_s_394;   // mult.v(1312)
    wire wfa_cout_394;   // mult.v(1312)
    wire wfa_s_395;   // mult.v(1313)
    wire wfa_cout_395;   // mult.v(1313)
    wire wfa_s_396;   // mult.v(1314)
    wire wfa_cout_396;   // mult.v(1314)
    wire wfa_s_397;   // mult.v(1315)
    wire wfa_cout_397;   // mult.v(1315)
    wire wfa_s_398;   // mult.v(1316)
    wire wfa_cout_398;   // mult.v(1316)
    wire wfa_s_399;   // mult.v(1317)
    wire wfa_cout_399;   // mult.v(1317)
    wire wfa_s_400;   // mult.v(1318)
    wire wfa_cout_400;   // mult.v(1318)
    wire wfa_s_401;   // mult.v(1319)
    wire wfa_cout_401;   // mult.v(1319)
    wire wfa_s_402;   // mult.v(1320)
    wire wfa_cout_402;   // mult.v(1320)
    wire wfa_s_403;   // mult.v(1321)
    wire wfa_cout_403;   // mult.v(1321)
    wire wfa_s_404;   // mult.v(1322)
    wire wfa_cout_404;   // mult.v(1322)
    wire wfa_s_405;   // mult.v(1323)
    wire wfa_cout_405;   // mult.v(1323)
    wire wfa_s_406;   // mult.v(1324)
    wire wfa_cout_406;   // mult.v(1324)
    wire wfa_s_407;   // mult.v(1325)
    wire wfa_cout_407;   // mult.v(1325)
    wire wfa_s_408;   // mult.v(1326)
    wire wfa_cout_408;   // mult.v(1326)
    wire wfa_s_409;   // mult.v(1327)
    wire wfa_cout_409;   // mult.v(1327)
    wire wfa_s_410;   // mult.v(1328)
    wire wfa_cout_410;   // mult.v(1328)
    wire wfa_s_411;   // mult.v(1329)
    wire wfa_cout_411;   // mult.v(1329)
    wire wfa_s_412;   // mult.v(1330)
    wire wfa_cout_412;   // mult.v(1330)
    wire wfa_s_413;   // mult.v(1331)
    wire wfa_cout_413;   // mult.v(1331)
    wire wfa_s_414;   // mult.v(1332)
    wire wfa_cout_414;   // mult.v(1332)
    wire wfa_s_415;   // mult.v(1333)
    wire wfa_cout_415;   // mult.v(1333)
    wire wfa_s_416;   // mult.v(1334)
    wire wfa_cout_416;   // mult.v(1334)
    wire wfa_s_417;   // mult.v(1335)
    wire wfa_cout_417;   // mult.v(1335)
    wire wfa_s_418;   // mult.v(1336)
    wire wfa_cout_418;   // mult.v(1336)
    wire wfa_s_419;   // mult.v(1337)
    wire wfa_cout_419;   // mult.v(1337)
    wire wfa_s_420;   // mult.v(1338)
    wire wfa_cout_420;   // mult.v(1338)
    wire wfa_s_421;   // mult.v(1339)
    wire wfa_cout_421;   // mult.v(1339)
    wire wfa_s_422;   // mult.v(1340)
    wire wfa_cout_422;   // mult.v(1340)
    wire wfa_s_423;   // mult.v(1341)
    wire wfa_cout_423;   // mult.v(1341)
    wire wfa_s_424;   // mult.v(1342)
    wire wfa_cout_424;   // mult.v(1342)
    wire wfa_s_425;   // mult.v(1343)
    wire wfa_cout_425;   // mult.v(1343)
    wire wfa_s_426;   // mult.v(1344)
    wire wfa_cout_426;   // mult.v(1344)
    wire wfa_s_427;   // mult.v(1345)
    wire wfa_cout_427;   // mult.v(1345)
    wire wfa_s_428;   // mult.v(1346)
    wire wfa_cout_428;   // mult.v(1346)
    wire wfa_s_429;   // mult.v(1347)
    wire wfa_cout_429;   // mult.v(1347)
    wire wfa_s_430;   // mult.v(1348)
    wire wfa_cout_430;   // mult.v(1348)
    wire wfa_s_431;   // mult.v(1349)
    wire wfa_cout_431;   // mult.v(1349)
    wire wfa_s_432;   // mult.v(1350)
    wire wfa_cout_432;   // mult.v(1350)
    wire wfa_s_433;   // mult.v(1351)
    wire wfa_cout_433;   // mult.v(1351)
    wire wfa_s_434;   // mult.v(1352)
    wire wfa_cout_434;   // mult.v(1352)
    wire wfa_s_435;   // mult.v(1353)
    wire wfa_cout_435;   // mult.v(1353)
    wire wfa_s_436;   // mult.v(1354)
    wire wfa_cout_436;   // mult.v(1354)
    wire wfa_s_437;   // mult.v(1355)
    wire wfa_cout_437;   // mult.v(1355)
    wire wfa_s_438;   // mult.v(1356)
    wire wfa_cout_438;   // mult.v(1356)
    wire wfa_s_439;   // mult.v(1357)
    wire wfa_cout_439;   // mult.v(1357)
    wire wfa_s_440;   // mult.v(1358)
    wire wfa_cout_440;   // mult.v(1358)
    wire wfa_s_441;   // mult.v(1359)
    wire wfa_cout_441;   // mult.v(1359)
    wire wfa_s_442;   // mult.v(1360)
    wire wfa_cout_442;   // mult.v(1360)
    wire wfa_s_443;   // mult.v(1361)
    wire wfa_cout_443;   // mult.v(1361)
    wire wfa_s_444;   // mult.v(1362)
    wire wfa_cout_444;   // mult.v(1362)
    wire wfa_s_445;   // mult.v(1363)
    wire wfa_cout_445;   // mult.v(1363)
    wire wfa_s_446;   // mult.v(1364)
    wire wfa_cout_446;   // mult.v(1364)
    wire wfa_s_447;   // mult.v(1365)
    wire wfa_cout_447;   // mult.v(1365)
    wire wfa_s_448;   // mult.v(1366)
    wire wfa_cout_448;   // mult.v(1366)
    wire wfa_s_449;   // mult.v(1367)
    wire wfa_cout_449;   // mult.v(1367)
    wire wfa_s_450;   // mult.v(1368)
    wire wfa_cout_450;   // mult.v(1368)
    wire wfa_s_451;   // mult.v(1369)
    wire wfa_cout_451;   // mult.v(1369)
    wire wfa_s_452;   // mult.v(1370)
    wire wfa_cout_452;   // mult.v(1370)
    wire wfa_s_453;   // mult.v(1371)
    wire wfa_cout_453;   // mult.v(1371)
    wire wfa_s_454;   // mult.v(1372)
    wire wfa_cout_454;   // mult.v(1372)
    wire wfa_s_455;   // mult.v(1373)
    wire wfa_cout_455;   // mult.v(1373)
    wire wfa_s_456;   // mult.v(1374)
    wire wfa_cout_456;   // mult.v(1374)
    wire wfa_s_457;   // mult.v(1375)
    wire wfa_cout_457;   // mult.v(1375)
    wire wfa_s_458;   // mult.v(1376)
    wire wfa_cout_458;   // mult.v(1376)
    wire wfa_s_459;   // mult.v(1377)
    wire wfa_cout_459;   // mult.v(1377)
    wire wfa_s_460;   // mult.v(1378)
    wire wfa_cout_460;   // mult.v(1378)
    wire wfa_s_461;   // mult.v(1379)
    wire wfa_cout_461;   // mult.v(1379)
    wire wfa_s_462;   // mult.v(1380)
    wire wfa_cout_462;   // mult.v(1380)
    wire wfa_s_463;   // mult.v(1381)
    wire wfa_cout_463;   // mult.v(1381)
    wire wfa_s_464;   // mult.v(1382)
    wire wfa_cout_464;   // mult.v(1382)
    wire wfa_s_465;   // mult.v(1383)
    wire wfa_cout_465;   // mult.v(1383)
    wire wfa_s_466;   // mult.v(1384)
    wire wfa_cout_466;   // mult.v(1384)
    wire wfa_s_467;   // mult.v(1385)
    wire wfa_cout_467;   // mult.v(1385)
    wire wfa_s_468;   // mult.v(1386)
    wire wfa_cout_468;   // mult.v(1386)
    wire wfa_s_469;   // mult.v(1387)
    wire wfa_cout_469;   // mult.v(1387)
    wire wfa_s_470;   // mult.v(1388)
    wire wfa_cout_470;   // mult.v(1388)
    wire wfa_s_471;   // mult.v(1389)
    wire wfa_cout_471;   // mult.v(1389)
    wire wfa_s_472;   // mult.v(1390)
    wire wfa_cout_472;   // mult.v(1390)
    wire wfa_s_473;   // mult.v(1391)
    wire wfa_cout_473;   // mult.v(1391)
    wire wfa_s_474;   // mult.v(1392)
    wire wfa_cout_474;   // mult.v(1392)
    wire wfa_s_475;   // mult.v(1393)
    wire wfa_cout_475;   // mult.v(1393)
    wire wfa_s_476;   // mult.v(1394)
    wire wfa_cout_476;   // mult.v(1394)
    wire wfa_s_477;   // mult.v(1395)
    wire wfa_cout_477;   // mult.v(1395)
    wire wfa_s_478;   // mult.v(1396)
    wire wfa_cout_478;   // mult.v(1396)
    wire wfa_s_479;   // mult.v(1397)
    wire wfa_cout_479;   // mult.v(1397)
    wire wfa_s_480;   // mult.v(1398)
    wire wfa_cout_480;   // mult.v(1398)
    wire wfa_s_481;   // mult.v(1399)
    wire wfa_cout_481;   // mult.v(1399)
    wire wfa_s_482;   // mult.v(1400)
    wire wfa_cout_482;   // mult.v(1400)
    wire wfa_s_483;   // mult.v(1401)
    wire wfa_cout_483;   // mult.v(1401)
    wire wfa_s_484;   // mult.v(1402)
    wire wfa_cout_484;   // mult.v(1402)
    wire wfa_s_485;   // mult.v(1403)
    wire wfa_cout_485;   // mult.v(1403)
    wire wfa_s_486;   // mult.v(1404)
    wire wfa_cout_486;   // mult.v(1404)
    wire wfa_s_487;   // mult.v(1405)
    wire wfa_cout_487;   // mult.v(1405)
    wire wfa_s_488;   // mult.v(1406)
    wire wfa_cout_488;   // mult.v(1406)
    wire wfa_s_489;   // mult.v(1407)
    wire wfa_cout_489;   // mult.v(1407)
    wire wfa_s_490;   // mult.v(1408)
    wire wfa_cout_490;   // mult.v(1408)
    wire wfa_s_491;   // mult.v(1409)
    wire wfa_cout_491;   // mult.v(1409)
    wire wfa_s_492;   // mult.v(1410)
    wire wfa_cout_492;   // mult.v(1410)
    wire wfa_s_493;   // mult.v(1411)
    wire wfa_cout_493;   // mult.v(1411)
    wire wfa_s_494;   // mult.v(1412)
    wire wfa_cout_494;   // mult.v(1412)
    wire wfa_s_495;   // mult.v(1413)
    wire wfa_cout_495;   // mult.v(1413)
    wire wfa_s_496;   // mult.v(1414)
    wire wfa_cout_496;   // mult.v(1414)
    wire wfa_s_497;   // mult.v(1415)
    wire wfa_cout_497;   // mult.v(1415)
    wire wand_976;   // mult.v(1416)
    wire wand_1007;   // mult.v(1417)
    wire wfa_s_498;   // mult.v(1418)
    wire wfa_cout_498;   // mult.v(1418)
    wire wfa_s_499;   // mult.v(1419)
    wire wfa_cout_499;   // mult.v(1419)
    wire wfa_s_500;   // mult.v(1420)
    wire wfa_cout_500;   // mult.v(1420)
    wire wfa_s_501;   // mult.v(1421)
    wire wfa_cout_501;   // mult.v(1421)
    wire wand_915;   // mult.v(1422)
    wire wand_946;   // mult.v(1423)
    wire wand_977;   // mult.v(1424)
    wire wfa_s_502;   // mult.v(1425)
    wire wfa_cout_502;   // mult.v(1425)
    wire wand_1008;   // mult.v(1426)
    wire wfa_s_503;   // mult.v(1427)
    wire wfa_cout_503;   // mult.v(1427)
    wire wfa_s_504;   // mult.v(1428)
    wire wfa_cout_504;   // mult.v(1428)
    wire wfa_s_505;   // mult.v(1429)
    wire wfa_cout_505;   // mult.v(1429)
    wire wand_854;   // mult.v(1430)
    wire wand_885;   // mult.v(1431)
    wire wand_916;   // mult.v(1432)
    wire wfa_s_506;   // mult.v(1433)
    wire wfa_cout_506;   // mult.v(1433)
    wire wand_947;   // mult.v(1434)
    wire wand_978;   // mult.v(1435)
    wire wand_1009;   // mult.v(1436)
    wire wfa_s_507;   // mult.v(1437)
    wire wfa_cout_507;   // mult.v(1437)
    wire wfa_s_508;   // mult.v(1438)
    wire wfa_cout_508;   // mult.v(1438)
    wire wfa_s_509;   // mult.v(1439)
    wire wfa_cout_509;   // mult.v(1439)
    wire wand_793;   // mult.v(1440)
    wire wand_824;   // mult.v(1441)
    wire wand_855;   // mult.v(1442)
    wire wfa_s_510;   // mult.v(1443)
    wire wfa_cout_510;   // mult.v(1443)
    wire wand_886;   // mult.v(1444)
    wire wand_917;   // mult.v(1445)
    wire wand_948;   // mult.v(1446)
    wire wfa_s_511;   // mult.v(1447)
    wire wfa_cout_511;   // mult.v(1447)
    wire wand_979;   // mult.v(1448)
    wire wand_1010;   // mult.v(1449)
    wire wfa_s_512;   // mult.v(1450)
    wire wfa_cout_512;   // mult.v(1450)
    wire wfa_s_513;   // mult.v(1451)
    wire wfa_cout_513;   // mult.v(1451)
    wire wand_732;   // mult.v(1452)
    wire wand_763;   // mult.v(1453)
    wire wand_794;   // mult.v(1454)
    wire wfa_s_514;   // mult.v(1455)
    wire wfa_cout_514;   // mult.v(1455)
    wire wand_825;   // mult.v(1456)
    wire wand_856;   // mult.v(1457)
    wire wand_887;   // mult.v(1458)
    wire wfa_s_515;   // mult.v(1459)
    wire wfa_cout_515;   // mult.v(1459)
    wire wand_918;   // mult.v(1460)
    wire wand_949;   // mult.v(1461)
    wire wand_980;   // mult.v(1462)
    wire wfa_s_516;   // mult.v(1463)
    wire wfa_cout_516;   // mult.v(1463)
    wire wand_1011;   // mult.v(1464)
    wire wfa_s_517;   // mult.v(1465)
    wire wfa_cout_517;   // mult.v(1465)
    wire wand_671;   // mult.v(1466)
    wire wand_702;   // mult.v(1467)
    wire wand_733;   // mult.v(1468)
    wire wfa_s_518;   // mult.v(1469)
    wire wfa_cout_518;   // mult.v(1469)
    wire wand_764;   // mult.v(1470)
    wire wand_795;   // mult.v(1471)
    wire wand_826;   // mult.v(1472)
    wire wfa_s_519;   // mult.v(1473)
    wire wfa_cout_519;   // mult.v(1473)
    wire wand_857;   // mult.v(1474)
    wire wand_888;   // mult.v(1475)
    wire wand_919;   // mult.v(1476)
    wire wfa_s_520;   // mult.v(1477)
    wire wfa_cout_520;   // mult.v(1477)
    wire wand_950;   // mult.v(1478)
    wire wand_981;   // mult.v(1479)
    wire wand_1012;   // mult.v(1480)
    wire wfa_s_521;   // mult.v(1481)
    wire wfa_cout_521;   // mult.v(1481)
    wire wand_703;   // mult.v(1482)
    wire wand_734;   // mult.v(1483)
    wire wand_765;   // mult.v(1484)
    wire wfa_s_522;   // mult.v(1485)
    wire wfa_cout_522;   // mult.v(1485)
    wire wand_796;   // mult.v(1486)
    wire wand_827;   // mult.v(1487)
    wire wand_858;   // mult.v(1488)
    wire wfa_s_523;   // mult.v(1489)
    wire wfa_cout_523;   // mult.v(1489)
    wire wand_889;   // mult.v(1490)
    wire wand_920;   // mult.v(1491)
    wire wand_951;   // mult.v(1492)
    wire wfa_s_524;   // mult.v(1493)
    wire wfa_cout_524;   // mult.v(1493)
    wire wand_735;   // mult.v(1494)
    wire wand_766;   // mult.v(1495)
    wire wand_797;   // mult.v(1496)
    wire wfa_s_525;   // mult.v(1497)
    wire wfa_cout_525;   // mult.v(1497)
    wire wand_828;   // mult.v(1498)
    wire wand_859;   // mult.v(1499)
    wire wand_890;   // mult.v(1500)
    wire wfa_s_526;   // mult.v(1501)
    wire wfa_cout_526;   // mult.v(1501)
    wire wand_767;   // mult.v(1502)
    wire wand_798;   // mult.v(1503)
    wire wand_829;   // mult.v(1504)
    wire wfa_s_527;   // mult.v(1505)
    wire wfa_cout_527;   // mult.v(1505)
    wire wand_6;   // mult.v(1506)
    wire wand_37;   // mult.v(1507)
    wire wha_s_24;   // mult.v(1508)
    wire wha_c_24;   // mult.v(1508)
    wire wand_7;   // mult.v(1509)
    wire wand_38;   // mult.v(1510)
    wire wand_69;   // mult.v(1511)
    wire wfa_s_528;   // mult.v(1512)
    wire wfa_cout_528;   // mult.v(1512)
    wire wand_100;   // mult.v(1513)
    wire wand_131;   // mult.v(1514)
    wire wha_s_25;   // mult.v(1515)
    wire wha_c_25;   // mult.v(1515)
    wire wand_8;   // mult.v(1516)
    wire wand_39;   // mult.v(1517)
    wire wand_70;   // mult.v(1518)
    wire wfa_s_529;   // mult.v(1519)
    wire wfa_cout_529;   // mult.v(1519)
    wire wand_101;   // mult.v(1520)
    wire wand_132;   // mult.v(1521)
    wire wand_163;   // mult.v(1522)
    wire wfa_s_530;   // mult.v(1523)
    wire wfa_cout_530;   // mult.v(1523)
    wire wand_194;   // mult.v(1524)
    wire wand_225;   // mult.v(1525)
    wire wha_s_26;   // mult.v(1526)
    wire wha_c_26;   // mult.v(1526)
    wire wand_71;   // mult.v(1527)
    wire wand_102;   // mult.v(1528)
    wire wand_133;   // mult.v(1529)
    wire wfa_s_531;   // mult.v(1530)
    wire wfa_cout_531;   // mult.v(1530)
    wire wand_164;   // mult.v(1531)
    wire wand_195;   // mult.v(1532)
    wire wand_226;   // mult.v(1533)
    wire wfa_s_532;   // mult.v(1534)
    wire wfa_cout_532;   // mult.v(1534)
    wire wand_257;   // mult.v(1535)
    wire wand_288;   // mult.v(1536)
    wire wfa_s_533;   // mult.v(1537)
    wire wfa_cout_533;   // mult.v(1537)
    wire wand_165;   // mult.v(1538)
    wire wand_196;   // mult.v(1539)
    wire wand_227;   // mult.v(1540)
    wire wfa_s_534;   // mult.v(1541)
    wire wfa_cout_534;   // mult.v(1541)
    wire wand_258;   // mult.v(1542)
    wire wand_289;   // mult.v(1543)
    wire wand_320;   // mult.v(1544)
    wire wfa_s_535;   // mult.v(1545)
    wire wfa_cout_535;   // mult.v(1545)
    wire wfa_s_536;   // mult.v(1546)
    wire wfa_cout_536;   // mult.v(1546)
    wire wand_259;   // mult.v(1547)
    wire wand_290;   // mult.v(1548)
    wire wand_321;   // mult.v(1549)
    wire wfa_s_537;   // mult.v(1550)
    wire wfa_cout_537;   // mult.v(1550)
    wire wand_352;   // mult.v(1551)
    wire wfa_s_538;   // mult.v(1552)
    wire wfa_cout_538;   // mult.v(1552)
    wire wfa_s_539;   // mult.v(1553)
    wire wfa_cout_539;   // mult.v(1553)
    wire wand_353;   // mult.v(1554)
    wire wand_384;   // mult.v(1555)
    wire wfa_s_540;   // mult.v(1556)
    wire wfa_cout_540;   // mult.v(1556)
    wire wfa_s_541;   // mult.v(1557)
    wire wfa_cout_541;   // mult.v(1557)
    wire wfa_s_542;   // mult.v(1558)
    wire wfa_cout_542;   // mult.v(1558)
    wire wfa_s_543;   // mult.v(1559)
    wire wfa_cout_543;   // mult.v(1559)
    wire wfa_s_544;   // mult.v(1560)
    wire wfa_cout_544;   // mult.v(1560)
    wire wfa_s_545;   // mult.v(1561)
    wire wfa_cout_545;   // mult.v(1561)
    wire wfa_s_546;   // mult.v(1562)
    wire wfa_cout_546;   // mult.v(1562)
    wire wfa_s_547;   // mult.v(1563)
    wire wfa_cout_547;   // mult.v(1563)
    wire wfa_s_548;   // mult.v(1564)
    wire wfa_cout_548;   // mult.v(1564)
    wire wfa_s_549;   // mult.v(1565)
    wire wfa_cout_549;   // mult.v(1565)
    wire wfa_s_550;   // mult.v(1566)
    wire wfa_cout_550;   // mult.v(1566)
    wire wfa_s_551;   // mult.v(1567)
    wire wfa_cout_551;   // mult.v(1567)
    wire wfa_s_552;   // mult.v(1568)
    wire wfa_cout_552;   // mult.v(1568)
    wire wfa_s_553;   // mult.v(1569)
    wire wfa_cout_553;   // mult.v(1569)
    wire wfa_s_554;   // mult.v(1570)
    wire wfa_cout_554;   // mult.v(1570)
    wire wfa_s_555;   // mult.v(1571)
    wire wfa_cout_555;   // mult.v(1571)
    wire wfa_s_556;   // mult.v(1572)
    wire wfa_cout_556;   // mult.v(1572)
    wire wfa_s_557;   // mult.v(1573)
    wire wfa_cout_557;   // mult.v(1573)
    wire wfa_s_558;   // mult.v(1574)
    wire wfa_cout_558;   // mult.v(1574)
    wire wfa_s_559;   // mult.v(1575)
    wire wfa_cout_559;   // mult.v(1575)
    wire wfa_s_560;   // mult.v(1576)
    wire wfa_cout_560;   // mult.v(1576)
    wire wfa_s_561;   // mult.v(1577)
    wire wfa_cout_561;   // mult.v(1577)
    wire wfa_s_562;   // mult.v(1578)
    wire wfa_cout_562;   // mult.v(1578)
    wire wfa_s_563;   // mult.v(1579)
    wire wfa_cout_563;   // mult.v(1579)
    wire wfa_s_564;   // mult.v(1580)
    wire wfa_cout_564;   // mult.v(1580)
    wire wfa_s_565;   // mult.v(1581)
    wire wfa_cout_565;   // mult.v(1581)
    wire wfa_s_566;   // mult.v(1582)
    wire wfa_cout_566;   // mult.v(1582)
    wire wfa_s_567;   // mult.v(1583)
    wire wfa_cout_567;   // mult.v(1583)
    wire wfa_s_568;   // mult.v(1584)
    wire wfa_cout_568;   // mult.v(1584)
    wire wfa_s_569;   // mult.v(1585)
    wire wfa_cout_569;   // mult.v(1585)
    wire wfa_s_570;   // mult.v(1586)
    wire wfa_cout_570;   // mult.v(1586)
    wire wfa_s_571;   // mult.v(1587)
    wire wfa_cout_571;   // mult.v(1587)
    wire wfa_s_572;   // mult.v(1588)
    wire wfa_cout_572;   // mult.v(1588)
    wire wfa_s_573;   // mult.v(1589)
    wire wfa_cout_573;   // mult.v(1589)
    wire wfa_s_574;   // mult.v(1590)
    wire wfa_cout_574;   // mult.v(1590)
    wire wfa_s_575;   // mult.v(1591)
    wire wfa_cout_575;   // mult.v(1591)
    wire wfa_s_576;   // mult.v(1592)
    wire wfa_cout_576;   // mult.v(1592)
    wire wfa_s_577;   // mult.v(1593)
    wire wfa_cout_577;   // mult.v(1593)
    wire wfa_s_578;   // mult.v(1594)
    wire wfa_cout_578;   // mult.v(1594)
    wire wfa_s_579;   // mult.v(1595)
    wire wfa_cout_579;   // mult.v(1595)
    wire wfa_s_580;   // mult.v(1596)
    wire wfa_cout_580;   // mult.v(1596)
    wire wfa_s_581;   // mult.v(1597)
    wire wfa_cout_581;   // mult.v(1597)
    wire wfa_s_582;   // mult.v(1598)
    wire wfa_cout_582;   // mult.v(1598)
    wire wfa_s_583;   // mult.v(1599)
    wire wfa_cout_583;   // mult.v(1599)
    wire wfa_s_584;   // mult.v(1600)
    wire wfa_cout_584;   // mult.v(1600)
    wire wfa_s_585;   // mult.v(1601)
    wire wfa_cout_585;   // mult.v(1601)
    wire wfa_s_586;   // mult.v(1602)
    wire wfa_cout_586;   // mult.v(1602)
    wire wfa_s_587;   // mult.v(1603)
    wire wfa_cout_587;   // mult.v(1603)
    wire wfa_s_588;   // mult.v(1604)
    wire wfa_cout_588;   // mult.v(1604)
    wire wfa_s_589;   // mult.v(1605)
    wire wfa_cout_589;   // mult.v(1605)
    wire wfa_s_590;   // mult.v(1606)
    wire wfa_cout_590;   // mult.v(1606)
    wire wfa_s_591;   // mult.v(1607)
    wire wfa_cout_591;   // mult.v(1607)
    wire wfa_s_592;   // mult.v(1608)
    wire wfa_cout_592;   // mult.v(1608)
    wire wfa_s_593;   // mult.v(1609)
    wire wfa_cout_593;   // mult.v(1609)
    wire wfa_s_594;   // mult.v(1610)
    wire wfa_cout_594;   // mult.v(1610)
    wire wfa_s_595;   // mult.v(1611)
    wire wfa_cout_595;   // mult.v(1611)
    wire wfa_s_596;   // mult.v(1612)
    wire wfa_cout_596;   // mult.v(1612)
    wire wfa_s_597;   // mult.v(1613)
    wire wfa_cout_597;   // mult.v(1613)
    wire wfa_s_598;   // mult.v(1614)
    wire wfa_cout_598;   // mult.v(1614)
    wire wfa_s_599;   // mult.v(1615)
    wire wfa_cout_599;   // mult.v(1615)
    wire wfa_s_600;   // mult.v(1616)
    wire wfa_cout_600;   // mult.v(1616)
    wire wfa_s_601;   // mult.v(1617)
    wire wfa_cout_601;   // mult.v(1617)
    wire wfa_s_602;   // mult.v(1618)
    wire wfa_cout_602;   // mult.v(1618)
    wire wfa_s_603;   // mult.v(1619)
    wire wfa_cout_603;   // mult.v(1619)
    wire wfa_s_604;   // mult.v(1620)
    wire wfa_cout_604;   // mult.v(1620)
    wire wfa_s_605;   // mult.v(1621)
    wire wfa_cout_605;   // mult.v(1621)
    wire wfa_s_606;   // mult.v(1622)
    wire wfa_cout_606;   // mult.v(1622)
    wire wfa_s_607;   // mult.v(1623)
    wire wfa_cout_607;   // mult.v(1623)
    wire wfa_s_608;   // mult.v(1624)
    wire wfa_cout_608;   // mult.v(1624)
    wire wfa_s_609;   // mult.v(1625)
    wire wfa_cout_609;   // mult.v(1625)
    wire wfa_s_610;   // mult.v(1626)
    wire wfa_cout_610;   // mult.v(1626)
    wire wfa_s_611;   // mult.v(1627)
    wire wfa_cout_611;   // mult.v(1627)
    wire wfa_s_612;   // mult.v(1628)
    wire wfa_cout_612;   // mult.v(1628)
    wire wfa_s_613;   // mult.v(1629)
    wire wfa_cout_613;   // mult.v(1629)
    wire wfa_s_614;   // mult.v(1630)
    wire wfa_cout_614;   // mult.v(1630)
    wire wfa_s_615;   // mult.v(1631)
    wire wfa_cout_615;   // mult.v(1631)
    wire wfa_s_616;   // mult.v(1632)
    wire wfa_cout_616;   // mult.v(1632)
    wire wfa_s_617;   // mult.v(1633)
    wire wfa_cout_617;   // mult.v(1633)
    wire wfa_s_618;   // mult.v(1634)
    wire wfa_cout_618;   // mult.v(1634)
    wire wfa_s_619;   // mult.v(1635)
    wire wfa_cout_619;   // mult.v(1635)
    wire wfa_s_620;   // mult.v(1636)
    wire wfa_cout_620;   // mult.v(1636)
    wire wfa_s_621;   // mult.v(1637)
    wire wfa_cout_621;   // mult.v(1637)
    wire wfa_s_622;   // mult.v(1638)
    wire wfa_cout_622;   // mult.v(1638)
    wire wfa_s_623;   // mult.v(1639)
    wire wfa_cout_623;   // mult.v(1639)
    wire wfa_s_624;   // mult.v(1640)
    wire wfa_cout_624;   // mult.v(1640)
    wire wfa_s_625;   // mult.v(1641)
    wire wfa_cout_625;   // mult.v(1641)
    wire wfa_s_626;   // mult.v(1642)
    wire wfa_cout_626;   // mult.v(1642)
    wire wfa_s_627;   // mult.v(1643)
    wire wfa_cout_627;   // mult.v(1643)
    wire wfa_s_628;   // mult.v(1644)
    wire wfa_cout_628;   // mult.v(1644)
    wire wfa_s_629;   // mult.v(1645)
    wire wfa_cout_629;   // mult.v(1645)
    wire wfa_s_630;   // mult.v(1646)
    wire wfa_cout_630;   // mult.v(1646)
    wire wfa_s_631;   // mult.v(1647)
    wire wfa_cout_631;   // mult.v(1647)
    wire wfa_s_632;   // mult.v(1648)
    wire wfa_cout_632;   // mult.v(1648)
    wire wfa_s_633;   // mult.v(1649)
    wire wfa_cout_633;   // mult.v(1649)
    wire wfa_s_634;   // mult.v(1650)
    wire wfa_cout_634;   // mult.v(1650)
    wire wfa_s_635;   // mult.v(1651)
    wire wfa_cout_635;   // mult.v(1651)
    wire wfa_s_636;   // mult.v(1652)
    wire wfa_cout_636;   // mult.v(1652)
    wire wfa_s_637;   // mult.v(1653)
    wire wfa_cout_637;   // mult.v(1653)
    wire wfa_s_638;   // mult.v(1654)
    wire wfa_cout_638;   // mult.v(1654)
    wire wfa_s_639;   // mult.v(1655)
    wire wfa_cout_639;   // mult.v(1655)
    wire wfa_s_640;   // mult.v(1656)
    wire wfa_cout_640;   // mult.v(1656)
    wire wfa_s_641;   // mult.v(1657)
    wire wfa_cout_641;   // mult.v(1657)
    wire wfa_s_642;   // mult.v(1658)
    wire wfa_cout_642;   // mult.v(1658)
    wire wfa_s_643;   // mult.v(1659)
    wire wfa_cout_643;   // mult.v(1659)
    wire wfa_s_644;   // mult.v(1660)
    wire wfa_cout_644;   // mult.v(1660)
    wire wfa_s_645;   // mult.v(1661)
    wire wfa_cout_645;   // mult.v(1661)
    wire wfa_s_646;   // mult.v(1662)
    wire wfa_cout_646;   // mult.v(1662)
    wire wfa_s_647;   // mult.v(1663)
    wire wfa_cout_647;   // mult.v(1663)
    wire wfa_s_648;   // mult.v(1664)
    wire wfa_cout_648;   // mult.v(1664)
    wire wfa_s_649;   // mult.v(1665)
    wire wfa_cout_649;   // mult.v(1665)
    wire wfa_s_650;   // mult.v(1666)
    wire wfa_cout_650;   // mult.v(1666)
    wire wfa_s_651;   // mult.v(1667)
    wire wfa_cout_651;   // mult.v(1667)
    wire wfa_s_652;   // mult.v(1668)
    wire wfa_cout_652;   // mult.v(1668)
    wire wfa_s_653;   // mult.v(1669)
    wire wfa_cout_653;   // mult.v(1669)
    wire wfa_s_654;   // mult.v(1670)
    wire wfa_cout_654;   // mult.v(1670)
    wire wfa_s_655;   // mult.v(1671)
    wire wfa_cout_655;   // mult.v(1671)
    wire wfa_s_656;   // mult.v(1672)
    wire wfa_cout_656;   // mult.v(1672)
    wire wfa_s_657;   // mult.v(1673)
    wire wfa_cout_657;   // mult.v(1673)
    wire wfa_s_658;   // mult.v(1674)
    wire wfa_cout_658;   // mult.v(1674)
    wire wfa_s_659;   // mult.v(1675)
    wire wfa_cout_659;   // mult.v(1675)
    wire wand_982;   // mult.v(1676)
    wire wand_1013;   // mult.v(1677)
    wire wfa_s_660;   // mult.v(1678)
    wire wfa_cout_660;   // mult.v(1678)
    wire wfa_s_661;   // mult.v(1679)
    wire wfa_cout_661;   // mult.v(1679)
    wire wfa_s_662;   // mult.v(1680)
    wire wfa_cout_662;   // mult.v(1680)
    wire wand_921;   // mult.v(1681)
    wire wand_952;   // mult.v(1682)
    wire wand_983;   // mult.v(1683)
    wire wfa_s_663;   // mult.v(1684)
    wire wfa_cout_663;   // mult.v(1684)
    wire wand_1014;   // mult.v(1685)
    wire wfa_s_664;   // mult.v(1686)
    wire wfa_cout_664;   // mult.v(1686)
    wire wfa_s_665;   // mult.v(1687)
    wire wfa_cout_665;   // mult.v(1687)
    wire wand_860;   // mult.v(1688)
    wire wand_891;   // mult.v(1689)
    wire wand_922;   // mult.v(1690)
    wire wfa_s_666;   // mult.v(1691)
    wire wfa_cout_666;   // mult.v(1691)
    wire wand_953;   // mult.v(1692)
    wire wand_984;   // mult.v(1693)
    wire wand_1015;   // mult.v(1694)
    wire wfa_s_667;   // mult.v(1695)
    wire wfa_cout_667;   // mult.v(1695)
    wire wfa_s_668;   // mult.v(1696)
    wire wfa_cout_668;   // mult.v(1696)
    wire wand_799;   // mult.v(1697)
    wire wand_830;   // mult.v(1698)
    wire wand_861;   // mult.v(1699)
    wire wfa_s_669;   // mult.v(1700)
    wire wfa_cout_669;   // mult.v(1700)
    wire wand_892;   // mult.v(1701)
    wire wand_923;   // mult.v(1702)
    wire wand_954;   // mult.v(1703)
    wire wfa_s_670;   // mult.v(1704)
    wire wfa_cout_670;   // mult.v(1704)
    wire wand_985;   // mult.v(1705)
    wire wand_1016;   // mult.v(1706)
    wire wfa_s_671;   // mult.v(1707)
    wire wfa_cout_671;   // mult.v(1707)
    wire wand_831;   // mult.v(1708)
    wire wand_862;   // mult.v(1709)
    wire wand_893;   // mult.v(1710)
    wire wfa_s_672;   // mult.v(1711)
    wire wfa_cout_672;   // mult.v(1711)
    wire wand_924;   // mult.v(1712)
    wire wand_955;   // mult.v(1713)
    wire wand_986;   // mult.v(1714)
    wire wfa_s_673;   // mult.v(1715)
    wire wfa_cout_673;   // mult.v(1715)
    wire wand_863;   // mult.v(1716)
    wire wand_894;   // mult.v(1717)
    wire wand_925;   // mult.v(1718)
    wire wfa_s_674;   // mult.v(1719)
    wire wfa_cout_674;   // mult.v(1719)
    wire wand_4;   // mult.v(1720)
    wire wand_35;   // mult.v(1721)
    wire wha_s_27;   // mult.v(1722)
    wire wha_c_27;   // mult.v(1722)
    wire wand_5;   // mult.v(1723)
    wire wand_36;   // mult.v(1724)
    wire wand_67;   // mult.v(1725)
    wire wfa_s_675;   // mult.v(1726)
    wire wfa_cout_675;   // mult.v(1726)
    wire wand_98;   // mult.v(1727)
    wire wand_129;   // mult.v(1728)
    wire wha_s_28;   // mult.v(1729)
    wire wha_c_28;   // mult.v(1729)
    wire wand_68;   // mult.v(1730)
    wire wand_99;   // mult.v(1731)
    wire wand_130;   // mult.v(1732)
    wire wfa_s_676;   // mult.v(1733)
    wire wfa_cout_676;   // mult.v(1733)
    wire wand_161;   // mult.v(1734)
    wire wand_192;   // mult.v(1735)
    wire wfa_s_677;   // mult.v(1736)
    wire wfa_cout_677;   // mult.v(1736)
    wire wand_162;   // mult.v(1737)
    wire wand_193;   // mult.v(1738)
    wire wand_224;   // mult.v(1739)
    wire wfa_s_678;   // mult.v(1740)
    wire wfa_cout_678;   // mult.v(1740)
    wire wfa_s_679;   // mult.v(1741)
    wire wfa_cout_679;   // mult.v(1741)
    wire wand_256;   // mult.v(1742)
    wire wfa_s_680;   // mult.v(1743)
    wire wfa_cout_680;   // mult.v(1743)
    wire wfa_s_681;   // mult.v(1744)
    wire wfa_cout_681;   // mult.v(1744)
    wire wfa_s_682;   // mult.v(1745)
    wire wfa_cout_682;   // mult.v(1745)
    wire wfa_s_683;   // mult.v(1746)
    wire wfa_cout_683;   // mult.v(1746)
    wire wfa_s_684;   // mult.v(1747)
    wire wfa_cout_684;   // mult.v(1747)
    wire wfa_s_685;   // mult.v(1748)
    wire wfa_cout_685;   // mult.v(1748)
    wire wfa_s_686;   // mult.v(1749)
    wire wfa_cout_686;   // mult.v(1749)
    wire wfa_s_687;   // mult.v(1750)
    wire wfa_cout_687;   // mult.v(1750)
    wire wfa_s_688;   // mult.v(1751)
    wire wfa_cout_688;   // mult.v(1751)
    wire wfa_s_689;   // mult.v(1752)
    wire wfa_cout_689;   // mult.v(1752)
    wire wfa_s_690;   // mult.v(1753)
    wire wfa_cout_690;   // mult.v(1753)
    wire wfa_s_691;   // mult.v(1754)
    wire wfa_cout_691;   // mult.v(1754)
    wire wfa_s_692;   // mult.v(1755)
    wire wfa_cout_692;   // mult.v(1755)
    wire wfa_s_693;   // mult.v(1756)
    wire wfa_cout_693;   // mult.v(1756)
    wire wfa_s_694;   // mult.v(1757)
    wire wfa_cout_694;   // mult.v(1757)
    wire wfa_s_695;   // mult.v(1758)
    wire wfa_cout_695;   // mult.v(1758)
    wire wfa_s_696;   // mult.v(1759)
    wire wfa_cout_696;   // mult.v(1759)
    wire wfa_s_697;   // mult.v(1760)
    wire wfa_cout_697;   // mult.v(1760)
    wire wfa_s_698;   // mult.v(1761)
    wire wfa_cout_698;   // mult.v(1761)
    wire wfa_s_699;   // mult.v(1762)
    wire wfa_cout_699;   // mult.v(1762)
    wire wfa_s_700;   // mult.v(1763)
    wire wfa_cout_700;   // mult.v(1763)
    wire wfa_s_701;   // mult.v(1764)
    wire wfa_cout_701;   // mult.v(1764)
    wire wfa_s_702;   // mult.v(1765)
    wire wfa_cout_702;   // mult.v(1765)
    wire wfa_s_703;   // mult.v(1766)
    wire wfa_cout_703;   // mult.v(1766)
    wire wfa_s_704;   // mult.v(1767)
    wire wfa_cout_704;   // mult.v(1767)
    wire wfa_s_705;   // mult.v(1768)
    wire wfa_cout_705;   // mult.v(1768)
    wire wfa_s_706;   // mult.v(1769)
    wire wfa_cout_706;   // mult.v(1769)
    wire wfa_s_707;   // mult.v(1770)
    wire wfa_cout_707;   // mult.v(1770)
    wire wfa_s_708;   // mult.v(1771)
    wire wfa_cout_708;   // mult.v(1771)
    wire wfa_s_709;   // mult.v(1772)
    wire wfa_cout_709;   // mult.v(1772)
    wire wfa_s_710;   // mult.v(1773)
    wire wfa_cout_710;   // mult.v(1773)
    wire wfa_s_711;   // mult.v(1774)
    wire wfa_cout_711;   // mult.v(1774)
    wire wfa_s_712;   // mult.v(1775)
    wire wfa_cout_712;   // mult.v(1775)
    wire wfa_s_713;   // mult.v(1776)
    wire wfa_cout_713;   // mult.v(1776)
    wire wfa_s_714;   // mult.v(1777)
    wire wfa_cout_714;   // mult.v(1777)
    wire wfa_s_715;   // mult.v(1778)
    wire wfa_cout_715;   // mult.v(1778)
    wire wfa_s_716;   // mult.v(1779)
    wire wfa_cout_716;   // mult.v(1779)
    wire wfa_s_717;   // mult.v(1780)
    wire wfa_cout_717;   // mult.v(1780)
    wire wfa_s_718;   // mult.v(1781)
    wire wfa_cout_718;   // mult.v(1781)
    wire wfa_s_719;   // mult.v(1782)
    wire wfa_cout_719;   // mult.v(1782)
    wire wfa_s_720;   // mult.v(1783)
    wire wfa_cout_720;   // mult.v(1783)
    wire wfa_s_721;   // mult.v(1784)
    wire wfa_cout_721;   // mult.v(1784)
    wire wfa_s_722;   // mult.v(1785)
    wire wfa_cout_722;   // mult.v(1785)
    wire wfa_s_723;   // mult.v(1786)
    wire wfa_cout_723;   // mult.v(1786)
    wire wfa_s_724;   // mult.v(1787)
    wire wfa_cout_724;   // mult.v(1787)
    wire wfa_s_725;   // mult.v(1788)
    wire wfa_cout_725;   // mult.v(1788)
    wire wfa_s_726;   // mult.v(1789)
    wire wfa_cout_726;   // mult.v(1789)
    wire wfa_s_727;   // mult.v(1790)
    wire wfa_cout_727;   // mult.v(1790)
    wire wfa_s_728;   // mult.v(1791)
    wire wfa_cout_728;   // mult.v(1791)
    wire wfa_s_729;   // mult.v(1792)
    wire wfa_cout_729;   // mult.v(1792)
    wire wfa_s_730;   // mult.v(1793)
    wire wfa_cout_730;   // mult.v(1793)
    wire wfa_s_731;   // mult.v(1794)
    wire wfa_cout_731;   // mult.v(1794)
    wire wfa_s_732;   // mult.v(1795)
    wire wfa_cout_732;   // mult.v(1795)
    wire wfa_s_733;   // mult.v(1796)
    wire wfa_cout_733;   // mult.v(1796)
    wire wfa_s_734;   // mult.v(1797)
    wire wfa_cout_734;   // mult.v(1797)
    wire wfa_s_735;   // mult.v(1798)
    wire wfa_cout_735;   // mult.v(1798)
    wire wfa_s_736;   // mult.v(1799)
    wire wfa_cout_736;   // mult.v(1799)
    wire wfa_s_737;   // mult.v(1800)
    wire wfa_cout_737;   // mult.v(1800)
    wire wfa_s_738;   // mult.v(1801)
    wire wfa_cout_738;   // mult.v(1801)
    wire wfa_s_739;   // mult.v(1802)
    wire wfa_cout_739;   // mult.v(1802)
    wire wfa_s_740;   // mult.v(1803)
    wire wfa_cout_740;   // mult.v(1803)
    wire wfa_s_741;   // mult.v(1804)
    wire wfa_cout_741;   // mult.v(1804)
    wire wfa_s_742;   // mult.v(1805)
    wire wfa_cout_742;   // mult.v(1805)
    wire wfa_s_743;   // mult.v(1806)
    wire wfa_cout_743;   // mult.v(1806)
    wire wfa_s_744;   // mult.v(1807)
    wire wfa_cout_744;   // mult.v(1807)
    wire wfa_s_745;   // mult.v(1808)
    wire wfa_cout_745;   // mult.v(1808)
    wire wfa_s_746;   // mult.v(1809)
    wire wfa_cout_746;   // mult.v(1809)
    wire wfa_s_747;   // mult.v(1810)
    wire wfa_cout_747;   // mult.v(1810)
    wire wfa_s_748;   // mult.v(1811)
    wire wfa_cout_748;   // mult.v(1811)
    wire wfa_s_749;   // mult.v(1812)
    wire wfa_cout_749;   // mult.v(1812)
    wire wfa_s_750;   // mult.v(1813)
    wire wfa_cout_750;   // mult.v(1813)
    wire wfa_s_751;   // mult.v(1814)
    wire wfa_cout_751;   // mult.v(1814)
    wire wfa_s_752;   // mult.v(1815)
    wire wfa_cout_752;   // mult.v(1815)
    wire wfa_s_753;   // mult.v(1816)
    wire wfa_cout_753;   // mult.v(1816)
    wire wfa_s_754;   // mult.v(1817)
    wire wfa_cout_754;   // mult.v(1817)
    wire wfa_s_755;   // mult.v(1818)
    wire wfa_cout_755;   // mult.v(1818)
    wire wfa_s_756;   // mult.v(1819)
    wire wfa_cout_756;   // mult.v(1819)
    wire wfa_s_757;   // mult.v(1820)
    wire wfa_cout_757;   // mult.v(1820)
    wire wfa_s_758;   // mult.v(1821)
    wire wfa_cout_758;   // mult.v(1821)
    wire wfa_s_759;   // mult.v(1822)
    wire wfa_cout_759;   // mult.v(1822)
    wire wfa_s_760;   // mult.v(1823)
    wire wfa_cout_760;   // mult.v(1823)
    wire wfa_s_761;   // mult.v(1824)
    wire wfa_cout_761;   // mult.v(1824)
    wire wfa_s_762;   // mult.v(1825)
    wire wfa_cout_762;   // mult.v(1825)
    wire wfa_s_763;   // mult.v(1826)
    wire wfa_cout_763;   // mult.v(1826)
    wire wfa_s_764;   // mult.v(1827)
    wire wfa_cout_764;   // mult.v(1827)
    wire wfa_s_765;   // mult.v(1828)
    wire wfa_cout_765;   // mult.v(1828)
    wire wfa_s_766;   // mult.v(1829)
    wire wfa_cout_766;   // mult.v(1829)
    wire wfa_s_767;   // mult.v(1830)
    wire wfa_cout_767;   // mult.v(1830)
    wire wfa_s_768;   // mult.v(1831)
    wire wfa_cout_768;   // mult.v(1831)
    wire wfa_s_769;   // mult.v(1832)
    wire wfa_cout_769;   // mult.v(1832)
    wire wfa_s_770;   // mult.v(1833)
    wire wfa_cout_770;   // mult.v(1833)
    wire wfa_s_771;   // mult.v(1834)
    wire wfa_cout_771;   // mult.v(1834)
    wire wfa_s_772;   // mult.v(1835)
    wire wfa_cout_772;   // mult.v(1835)
    wire wfa_s_773;   // mult.v(1836)
    wire wfa_cout_773;   // mult.v(1836)
    wire wfa_s_774;   // mult.v(1837)
    wire wfa_cout_774;   // mult.v(1837)
    wire wfa_s_775;   // mult.v(1838)
    wire wfa_cout_775;   // mult.v(1838)
    wire wand_1017;   // mult.v(1839)
    wire wfa_s_776;   // mult.v(1840)
    wire wfa_cout_776;   // mult.v(1840)
    wire wfa_s_777;   // mult.v(1841)
    wire wfa_cout_777;   // mult.v(1841)
    wire wand_956;   // mult.v(1842)
    wire wand_987;   // mult.v(1843)
    wire wand_1018;   // mult.v(1844)
    wire wfa_s_778;   // mult.v(1845)
    wire wfa_cout_778;   // mult.v(1845)
    wire wfa_s_779;   // mult.v(1846)
    wire wfa_cout_779;   // mult.v(1846)
    wire wand_895;   // mult.v(1847)
    wire wand_926;   // mult.v(1848)
    wire wand_957;   // mult.v(1849)
    wire wfa_s_780;   // mult.v(1850)
    wire wfa_cout_780;   // mult.v(1850)
    wire wand_988;   // mult.v(1851)
    wire wand_1019;   // mult.v(1852)
    wire wfa_s_781;   // mult.v(1853)
    wire wfa_cout_781;   // mult.v(1853)
    wire wand_927;   // mult.v(1854)
    wire wand_958;   // mult.v(1855)
    wire wand_989;   // mult.v(1856)
    wire wfa_s_782;   // mult.v(1857)
    wire wfa_cout_782;   // mult.v(1857)
    wire wand_3;   // mult.v(1858)
    wire wand_34;   // mult.v(1859)
    wire wha_s_29;   // mult.v(1860)
    wire wha_c_29;   // mult.v(1860)
    wire wand_66;   // mult.v(1861)
    wire wand_97;   // mult.v(1862)
    wire wand_128;   // mult.v(1863)
    wire wfa_s_783;   // mult.v(1864)
    wire wfa_cout_783;   // mult.v(1864)
    wire wand_160;   // mult.v(1865)
    wire wfa_s_784;   // mult.v(1866)
    wire wfa_cout_784;   // mult.v(1866)
    wire wfa_s_785;   // mult.v(1867)
    wire wfa_cout_785;   // mult.v(1867)
    wire wfa_s_786;   // mult.v(1868)
    wire wfa_cout_786;   // mult.v(1868)
    wire wfa_s_787;   // mult.v(1869)
    wire wfa_cout_787;   // mult.v(1869)
    wire wfa_s_788;   // mult.v(1870)
    wire wfa_cout_788;   // mult.v(1870)
    wire wfa_s_789;   // mult.v(1871)
    wire wfa_cout_789;   // mult.v(1871)
    wire wfa_s_790;   // mult.v(1872)
    wire wfa_cout_790;   // mult.v(1872)
    wire wfa_s_791;   // mult.v(1873)
    wire wfa_cout_791;   // mult.v(1873)
    wire wfa_s_792;   // mult.v(1874)
    wire wfa_cout_792;   // mult.v(1874)
    wire wfa_s_793;   // mult.v(1875)
    wire wfa_cout_793;   // mult.v(1875)
    wire wfa_s_794;   // mult.v(1876)
    wire wfa_cout_794;   // mult.v(1876)
    wire wfa_s_795;   // mult.v(1877)
    wire wfa_cout_795;   // mult.v(1877)
    wire wfa_s_796;   // mult.v(1878)
    wire wfa_cout_796;   // mult.v(1878)
    wire wfa_s_797;   // mult.v(1879)
    wire wfa_cout_797;   // mult.v(1879)
    wire wfa_s_798;   // mult.v(1880)
    wire wfa_cout_798;   // mult.v(1880)
    wire wfa_s_799;   // mult.v(1881)
    wire wfa_cout_799;   // mult.v(1881)
    wire wfa_s_800;   // mult.v(1882)
    wire wfa_cout_800;   // mult.v(1882)
    wire wfa_s_801;   // mult.v(1883)
    wire wfa_cout_801;   // mult.v(1883)
    wire wfa_s_802;   // mult.v(1884)
    wire wfa_cout_802;   // mult.v(1884)
    wire wfa_s_803;   // mult.v(1885)
    wire wfa_cout_803;   // mult.v(1885)
    wire wfa_s_804;   // mult.v(1886)
    wire wfa_cout_804;   // mult.v(1886)
    wire wfa_s_805;   // mult.v(1887)
    wire wfa_cout_805;   // mult.v(1887)
    wire wfa_s_806;   // mult.v(1888)
    wire wfa_cout_806;   // mult.v(1888)
    wire wfa_s_807;   // mult.v(1889)
    wire wfa_cout_807;   // mult.v(1889)
    wire wfa_s_808;   // mult.v(1890)
    wire wfa_cout_808;   // mult.v(1890)
    wire wfa_s_809;   // mult.v(1891)
    wire wfa_cout_809;   // mult.v(1891)
    wire wfa_s_810;   // mult.v(1892)
    wire wfa_cout_810;   // mult.v(1892)
    wire wfa_s_811;   // mult.v(1893)
    wire wfa_cout_811;   // mult.v(1893)
    wire wfa_s_812;   // mult.v(1894)
    wire wfa_cout_812;   // mult.v(1894)
    wire wfa_s_813;   // mult.v(1895)
    wire wfa_cout_813;   // mult.v(1895)
    wire wfa_s_814;   // mult.v(1896)
    wire wfa_cout_814;   // mult.v(1896)
    wire wfa_s_815;   // mult.v(1897)
    wire wfa_cout_815;   // mult.v(1897)
    wire wfa_s_816;   // mult.v(1898)
    wire wfa_cout_816;   // mult.v(1898)
    wire wfa_s_817;   // mult.v(1899)
    wire wfa_cout_817;   // mult.v(1899)
    wire wfa_s_818;   // mult.v(1900)
    wire wfa_cout_818;   // mult.v(1900)
    wire wfa_s_819;   // mult.v(1901)
    wire wfa_cout_819;   // mult.v(1901)
    wire wfa_s_820;   // mult.v(1902)
    wire wfa_cout_820;   // mult.v(1902)
    wire wfa_s_821;   // mult.v(1903)
    wire wfa_cout_821;   // mult.v(1903)
    wire wfa_s_822;   // mult.v(1904)
    wire wfa_cout_822;   // mult.v(1904)
    wire wfa_s_823;   // mult.v(1905)
    wire wfa_cout_823;   // mult.v(1905)
    wire wfa_s_824;   // mult.v(1906)
    wire wfa_cout_824;   // mult.v(1906)
    wire wfa_s_825;   // mult.v(1907)
    wire wfa_cout_825;   // mult.v(1907)
    wire wfa_s_826;   // mult.v(1908)
    wire wfa_cout_826;   // mult.v(1908)
    wire wfa_s_827;   // mult.v(1909)
    wire wfa_cout_827;   // mult.v(1909)
    wire wfa_s_828;   // mult.v(1910)
    wire wfa_cout_828;   // mult.v(1910)
    wire wfa_s_829;   // mult.v(1911)
    wire wfa_cout_829;   // mult.v(1911)
    wire wfa_s_830;   // mult.v(1912)
    wire wfa_cout_830;   // mult.v(1912)
    wire wfa_s_831;   // mult.v(1913)
    wire wfa_cout_831;   // mult.v(1913)
    wire wfa_s_832;   // mult.v(1914)
    wire wfa_cout_832;   // mult.v(1914)
    wire wfa_s_833;   // mult.v(1915)
    wire wfa_cout_833;   // mult.v(1915)
    wire wfa_s_834;   // mult.v(1916)
    wire wfa_cout_834;   // mult.v(1916)
    wire wfa_s_835;   // mult.v(1917)
    wire wfa_cout_835;   // mult.v(1917)
    wire wfa_s_836;   // mult.v(1918)
    wire wfa_cout_836;   // mult.v(1918)
    wire wfa_s_837;   // mult.v(1919)
    wire wfa_cout_837;   // mult.v(1919)
    wire wand_1020;   // mult.v(1920)
    wire wfa_s_838;   // mult.v(1921)
    wire wfa_cout_838;   // mult.v(1921)
    wire wand_959;   // mult.v(1922)
    wire wand_990;   // mult.v(1923)
    wire wand_1021;   // mult.v(1924)
    wire wfa_s_839;   // mult.v(1925)
    wire wfa_cout_839;   // mult.v(1925)
    wire wand_2;   // mult.v(1926)
    wire wand_33;   // mult.v(1927)
    wire wha_s_30;   // mult.v(1928)
    wire wha_c_30;   // mult.v(1928)
    wire wand_65;   // mult.v(1929)
    wire wand_96;   // mult.v(1930)
    wire wfa_s_840;   // mult.v(1931)
    wire wfa_cout_840;   // mult.v(1931)
    wire wfa_s_841;   // mult.v(1932)
    wire wfa_cout_841;   // mult.v(1932)
    wire wfa_s_842;   // mult.v(1933)
    wire wfa_cout_842;   // mult.v(1933)
    wire wfa_s_843;   // mult.v(1934)
    wire wfa_cout_843;   // mult.v(1934)
    wire wfa_s_844;   // mult.v(1935)
    wire wfa_cout_844;   // mult.v(1935)
    wire wfa_s_845;   // mult.v(1936)
    wire wfa_cout_845;   // mult.v(1936)
    wire wfa_s_846;   // mult.v(1937)
    wire wfa_cout_846;   // mult.v(1937)
    wire wfa_s_847;   // mult.v(1938)
    wire wfa_cout_847;   // mult.v(1938)
    wire wfa_s_848;   // mult.v(1939)
    wire wfa_cout_848;   // mult.v(1939)
    wire wfa_s_849;   // mult.v(1940)
    wire wfa_cout_849;   // mult.v(1940)
    wire wfa_s_850;   // mult.v(1941)
    wire wfa_cout_850;   // mult.v(1941)
    wire wfa_s_851;   // mult.v(1942)
    wire wfa_cout_851;   // mult.v(1942)
    wire wfa_s_852;   // mult.v(1943)
    wire wfa_cout_852;   // mult.v(1943)
    wire wfa_s_853;   // mult.v(1944)
    wire wfa_cout_853;   // mult.v(1944)
    wire wfa_s_854;   // mult.v(1945)
    wire wfa_cout_854;   // mult.v(1945)
    wire wfa_s_855;   // mult.v(1946)
    wire wfa_cout_855;   // mult.v(1946)
    wire wfa_s_856;   // mult.v(1947)
    wire wfa_cout_856;   // mult.v(1947)
    wire wfa_s_857;   // mult.v(1948)
    wire wfa_cout_857;   // mult.v(1948)
    wire wfa_s_858;   // mult.v(1949)
    wire wfa_cout_858;   // mult.v(1949)
    wire wfa_s_859;   // mult.v(1950)
    wire wfa_cout_859;   // mult.v(1950)
    wire wfa_s_860;   // mult.v(1951)
    wire wfa_cout_860;   // mult.v(1951)
    wire wfa_s_861;   // mult.v(1952)
    wire wfa_cout_861;   // mult.v(1952)
    wire wfa_s_862;   // mult.v(1953)
    wire wfa_cout_862;   // mult.v(1953)
    wire wfa_s_863;   // mult.v(1954)
    wire wfa_cout_863;   // mult.v(1954)
    wire wfa_s_864;   // mult.v(1955)
    wire wfa_cout_864;   // mult.v(1955)
    wire wfa_s_865;   // mult.v(1956)
    wire wfa_cout_865;   // mult.v(1956)
    wire wfa_s_866;   // mult.v(1957)
    wire wfa_cout_866;   // mult.v(1957)
    wire wfa_s_867;   // mult.v(1958)
    wire wfa_cout_867;   // mult.v(1958)
    wire wfa_s_868;   // mult.v(1959)
    wire wfa_cout_868;   // mult.v(1959)
    wire wfa_s_869;   // mult.v(1960)
    wire wfa_cout_869;   // mult.v(1960)
    wire wfa_s_870;   // mult.v(1961)
    wire wfa_cout_870;   // mult.v(1961)
    wire wfa_s_871;   // mult.v(1962)
    wire wfa_cout_871;   // mult.v(1962)
    wire wfa_s_872;   // mult.v(1963)
    wire wfa_cout_872;   // mult.v(1963)
    wire wfa_s_873;   // mult.v(1964)
    wire wfa_cout_873;   // mult.v(1964)
    wire wfa_s_874;   // mult.v(1965)
    wire wfa_cout_874;   // mult.v(1965)
    wire wfa_s_875;   // mult.v(1966)
    wire wfa_cout_875;   // mult.v(1966)
    wire wfa_s_876;   // mult.v(1967)
    wire wfa_cout_876;   // mult.v(1967)
    wire wfa_s_877;   // mult.v(1968)
    wire wfa_cout_877;   // mult.v(1968)
    wire wfa_s_878;   // mult.v(1969)
    wire wfa_cout_878;   // mult.v(1969)
    wire wfa_s_879;   // mult.v(1970)
    wire wfa_cout_879;   // mult.v(1970)
    wire wfa_s_880;   // mult.v(1971)
    wire wfa_cout_880;   // mult.v(1971)
    wire wfa_s_881;   // mult.v(1972)
    wire wfa_cout_881;   // mult.v(1972)
    wire wfa_s_882;   // mult.v(1973)
    wire wfa_cout_882;   // mult.v(1973)
    wire wfa_s_883;   // mult.v(1974)
    wire wfa_cout_883;   // mult.v(1974)
    wire wfa_s_884;   // mult.v(1975)
    wire wfa_cout_884;   // mult.v(1975)
    wire wfa_s_885;   // mult.v(1976)
    wire wfa_cout_885;   // mult.v(1976)
    wire wfa_s_886;   // mult.v(1977)
    wire wfa_cout_886;   // mult.v(1977)
    wire wfa_s_887;   // mult.v(1978)
    wire wfa_cout_887;   // mult.v(1978)
    wire wfa_s_888;   // mult.v(1979)
    wire wfa_cout_888;   // mult.v(1979)
    wire wfa_s_889;   // mult.v(1980)
    wire wfa_cout_889;   // mult.v(1980)
    wire wfa_s_890;   // mult.v(1981)
    wire wfa_cout_890;   // mult.v(1981)
    wire wfa_s_891;   // mult.v(1982)
    wire wfa_cout_891;   // mult.v(1982)
    wire wfa_s_892;   // mult.v(1983)
    wire wfa_cout_892;   // mult.v(1983)
    wire wfa_s_893;   // mult.v(1984)
    wire wfa_cout_893;   // mult.v(1984)
    wire wfa_s_894;   // mult.v(1985)
    wire wfa_cout_894;   // mult.v(1985)
    wire wfa_s_895;   // mult.v(1986)
    wire wfa_cout_895;   // mult.v(1986)
    wire wfa_s_896;   // mult.v(1987)
    wire wfa_cout_896;   // mult.v(1987)
    wire wfa_s_897;   // mult.v(1988)
    wire wfa_cout_897;   // mult.v(1988)
    wire wand_991;   // mult.v(1989)
    wire wand_1022;   // mult.v(1990)
    wire wfa_s_898;   // mult.v(1991)
    wire wfa_cout_898;   // mult.v(1991)
    wire wand_1;   // mult.v(1992)
    wire wand_32;   // mult.v(1993)
    wire wha_c_31;   // mult.v(1994)
    wire wand_64;   // mult.v(1995)
    wire wfa_cout_899;   // mult.v(1996)
    wire wfa_cout_900;   // mult.v(1997)
    wire wfa_cout_901;   // mult.v(1998)
    wire wfa_cout_902;   // mult.v(1999)
    wire wfa_cout_903;   // mult.v(2000)
    wire wfa_cout_904;   // mult.v(2001)
    wire wfa_cout_905;   // mult.v(2002)
    wire wfa_cout_906;   // mult.v(2003)
    wire wfa_cout_907;   // mult.v(2004)
    wire wfa_cout_908;   // mult.v(2005)
    wire wfa_cout_909;   // mult.v(2006)
    wire wfa_cout_910;   // mult.v(2007)
    wire wfa_cout_911;   // mult.v(2008)
    wire wfa_cout_912;   // mult.v(2009)
    wire wfa_cout_913;   // mult.v(2010)
    wire wfa_cout_914;   // mult.v(2011)
    wire wfa_cout_915;   // mult.v(2012)
    wire wfa_cout_916;   // mult.v(2013)
    wire wfa_cout_917;   // mult.v(2014)
    wire wfa_cout_918;   // mult.v(2015)
    wire wfa_cout_919;   // mult.v(2016)
    wire wfa_cout_920;   // mult.v(2017)
    wire wfa_cout_921;   // mult.v(2018)
    wire wfa_cout_922;   // mult.v(2019)
    wire wfa_cout_923;   // mult.v(2020)
    wire wfa_cout_924;   // mult.v(2021)
    wire wfa_cout_925;   // mult.v(2022)
    wire wfa_cout_926;   // mult.v(2023)
    wire wfa_cout_927;   // mult.v(2024)
    wire wfa_cout_928;   // mult.v(2025)
    wire wfa_cout_929;   // mult.v(2026)
    wire wfa_cout_930;   // mult.v(2027)
    wire wfa_cout_931;   // mult.v(2028)
    wire wfa_cout_932;   // mult.v(2029)
    wire wfa_cout_933;   // mult.v(2030)
    wire wfa_cout_934;   // mult.v(2031)
    wire wfa_cout_935;   // mult.v(2032)
    wire wfa_cout_936;   // mult.v(2033)
    wire wfa_cout_937;   // mult.v(2034)
    wire wfa_cout_938;   // mult.v(2035)
    wire wfa_cout_939;   // mult.v(2036)
    wire wfa_cout_940;   // mult.v(2037)
    wire wfa_cout_941;   // mult.v(2038)
    wire wfa_cout_942;   // mult.v(2039)
    wire wfa_cout_943;   // mult.v(2040)
    wire wfa_cout_944;   // mult.v(2041)
    wire wfa_cout_945;   // mult.v(2042)
    wire wfa_cout_946;   // mult.v(2043)
    wire wfa_cout_947;   // mult.v(2044)
    wire wfa_cout_948;   // mult.v(2045)
    wire wfa_cout_949;   // mult.v(2046)
    wire wfa_cout_950;   // mult.v(2047)
    wire wfa_cout_951;   // mult.v(2048)
    wire wfa_cout_952;   // mult.v(2049)
    wire wfa_cout_953;   // mult.v(2050)
    wire wfa_cout_954;   // mult.v(2051)
    wire wfa_cout_955;   // mult.v(2052)
    wire wfa_cout_956;   // mult.v(2053)
    wire wfa_cout_957;   // mult.v(2054)
    wire wfa_cout_958;   // mult.v(2055)
    wire wand_1023;   // mult.v(2056)
    
    and (wand_28, a[0], b[28]) ;   // mult.v(2060)
    and (wand_59, a[1], b[27]) ;   // mult.v(2061)
    ha ha_0 (.a(wand_28), .b(wand_59), .s(wha_s_0), .c(wha_c_0));   // mult.v(2062)
    and (wand_29, a[0], b[29]) ;   // mult.v(2063)
    and (wand_60, a[1], b[28]) ;   // mult.v(2064)
    and (wand_91, a[2], b[27]) ;   // mult.v(2065)
    fa fa_0 (.a(wand_29), .b(wand_60), .cin(wand_91), .s(wfa_s_0), .cout(wfa_cout_0));   // mult.v(2066)
    and (wand_122, a[3], b[26]) ;   // mult.v(2067)
    and (wand_153, a[4], b[25]) ;   // mult.v(2068)
    ha ha_1 (.a(wand_122), .b(wand_153), .s(wha_s_1), .c(wha_c_1));   // mult.v(2069)
    and (wand_30, a[0], b[30]) ;   // mult.v(2070)
    and (wand_61, a[1], b[29]) ;   // mult.v(2071)
    and (wand_92, a[2], b[28]) ;   // mult.v(2072)
    fa fa_1 (.a(wand_30), .b(wand_61), .cin(wand_92), .s(wfa_s_1), .cout(wfa_cout_1));   // mult.v(2073)
    and (wand_123, a[3], b[27]) ;   // mult.v(2074)
    and (wand_154, a[4], b[26]) ;   // mult.v(2075)
    and (wand_185, a[5], b[25]) ;   // mult.v(2076)
    fa fa_2 (.a(wand_123), .b(wand_154), .cin(wand_185), .s(wfa_s_2), 
       .cout(wfa_cout_2));   // mult.v(2077)
    and (wand_216, a[6], b[24]) ;   // mult.v(2078)
    and (wand_247, a[7], b[23]) ;   // mult.v(2079)
    ha ha_2 (.a(wand_216), .b(wand_247), .s(wha_s_2), .c(wha_c_2));   // mult.v(2080)
    and (wand_31, a[0], b[31]) ;   // mult.v(2081)
    and (wand_62, a[1], b[30]) ;   // mult.v(2082)
    and (wand_93, a[2], b[29]) ;   // mult.v(2083)
    fa fa_3 (.a(wand_31), .b(wand_62), .cin(wand_93), .s(wfa_s_3), .cout(wfa_cout_3));   // mult.v(2084)
    and (wand_124, a[3], b[28]) ;   // mult.v(2085)
    and (wand_155, a[4], b[27]) ;   // mult.v(2086)
    and (wand_186, a[5], b[26]) ;   // mult.v(2087)
    fa fa_4 (.a(wand_124), .b(wand_155), .cin(wand_186), .s(wfa_s_4), 
       .cout(wfa_cout_4));   // mult.v(2088)
    and (wand_217, a[6], b[25]) ;   // mult.v(2089)
    and (wand_248, a[7], b[24]) ;   // mult.v(2090)
    and (wand_279, a[8], b[23]) ;   // mult.v(2091)
    fa fa_5 (.a(wand_217), .b(wand_248), .cin(wand_279), .s(wfa_s_5), 
       .cout(wfa_cout_5));   // mult.v(2092)
    and (wand_310, a[9], b[22]) ;   // mult.v(2093)
    and (wand_341, a[10], b[21]) ;   // mult.v(2094)
    ha ha_3 (.a(wand_310), .b(wand_341), .s(wha_s_3), .c(wha_c_3));   // mult.v(2095)
    and (wand_63, a[1], b[31]) ;   // mult.v(2096)
    and (wand_94, a[2], b[30]) ;   // mult.v(2097)
    and (wand_125, a[3], b[29]) ;   // mult.v(2098)
    fa fa_6 (.a(wand_63), .b(wand_94), .cin(wand_125), .s(wfa_s_6), 
       .cout(wfa_cout_6));   // mult.v(2099)
    and (wand_156, a[4], b[28]) ;   // mult.v(2100)
    and (wand_187, a[5], b[27]) ;   // mult.v(2101)
    and (wand_218, a[6], b[26]) ;   // mult.v(2102)
    fa fa_7 (.a(wand_156), .b(wand_187), .cin(wand_218), .s(wfa_s_7), 
       .cout(wfa_cout_7));   // mult.v(2103)
    and (wand_249, a[7], b[25]) ;   // mult.v(2104)
    and (wand_280, a[8], b[24]) ;   // mult.v(2105)
    and (wand_311, a[9], b[23]) ;   // mult.v(2106)
    fa fa_8 (.a(wand_249), .b(wand_280), .cin(wand_311), .s(wfa_s_8), 
       .cout(wfa_cout_8));   // mult.v(2107)
    and (wand_342, a[10], b[22]) ;   // mult.v(2108)
    and (wand_373, a[11], b[21]) ;   // mult.v(2109)
    ha ha_4 (.a(wand_342), .b(wand_373), .s(wha_s_4), .c(wha_c_4));   // mult.v(2110)
    and (wand_95, a[2], b[31]) ;   // mult.v(2111)
    and (wand_126, a[3], b[30]) ;   // mult.v(2112)
    and (wand_157, a[4], b[29]) ;   // mult.v(2113)
    fa fa_9 (.a(wand_95), .b(wand_126), .cin(wand_157), .s(wfa_s_9), 
       .cout(wfa_cout_9));   // mult.v(2114)
    and (wand_188, a[5], b[28]) ;   // mult.v(2115)
    and (wand_219, a[6], b[27]) ;   // mult.v(2116)
    and (wand_250, a[7], b[26]) ;   // mult.v(2117)
    fa fa_10 (.a(wand_188), .b(wand_219), .cin(wand_250), .s(wfa_s_10), 
       .cout(wfa_cout_10));   // mult.v(2118)
    and (wand_281, a[8], b[25]) ;   // mult.v(2119)
    and (wand_312, a[9], b[24]) ;   // mult.v(2120)
    and (wand_343, a[10], b[23]) ;   // mult.v(2121)
    fa fa_11 (.a(wand_281), .b(wand_312), .cin(wand_343), .s(wfa_s_11), 
       .cout(wfa_cout_11));   // mult.v(2122)
    and (wand_127, a[3], b[31]) ;   // mult.v(2123)
    and (wand_158, a[4], b[30]) ;   // mult.v(2124)
    and (wand_189, a[5], b[29]) ;   // mult.v(2125)
    fa fa_12 (.a(wand_127), .b(wand_158), .cin(wand_189), .s(wfa_s_12), 
       .cout(wfa_cout_12));   // mult.v(2126)
    and (wand_220, a[6], b[28]) ;   // mult.v(2127)
    and (wand_251, a[7], b[27]) ;   // mult.v(2128)
    and (wand_282, a[8], b[26]) ;   // mult.v(2129)
    fa fa_13 (.a(wand_220), .b(wand_251), .cin(wand_282), .s(wfa_s_13), 
       .cout(wfa_cout_13));   // mult.v(2130)
    and (wand_159, a[4], b[31]) ;   // mult.v(2131)
    and (wand_190, a[5], b[30]) ;   // mult.v(2132)
    and (wand_221, a[6], b[29]) ;   // mult.v(2133)
    fa fa_14 (.a(wand_159), .b(wand_190), .cin(wand_221), .s(wfa_s_14), 
       .cout(wfa_cout_14));   // mult.v(2134)
    and (wand_19, a[0], b[19]) ;   // mult.v(2135)
    and (wand_50, a[1], b[18]) ;   // mult.v(2136)
    ha ha_5 (.a(wand_19), .b(wand_50), .s(wha_s_5), .c(wha_c_5));   // mult.v(2137)
    and (wand_20, a[0], b[20]) ;   // mult.v(2138)
    and (wand_51, a[1], b[19]) ;   // mult.v(2139)
    and (wand_82, a[2], b[18]) ;   // mult.v(2140)
    fa fa_15 (.a(wand_20), .b(wand_51), .cin(wand_82), .s(wfa_s_15), 
       .cout(wfa_cout_15));   // mult.v(2141)
    and (wand_113, a[3], b[17]) ;   // mult.v(2142)
    and (wand_144, a[4], b[16]) ;   // mult.v(2143)
    ha ha_6 (.a(wand_113), .b(wand_144), .s(wha_s_6), .c(wha_c_6));   // mult.v(2144)
    and (wand_21, a[0], b[21]) ;   // mult.v(2145)
    and (wand_52, a[1], b[20]) ;   // mult.v(2146)
    and (wand_83, a[2], b[19]) ;   // mult.v(2147)
    fa fa_16 (.a(wand_21), .b(wand_52), .cin(wand_83), .s(wfa_s_16), 
       .cout(wfa_cout_16));   // mult.v(2148)
    and (wand_114, a[3], b[18]) ;   // mult.v(2149)
    and (wand_145, a[4], b[17]) ;   // mult.v(2150)
    and (wand_176, a[5], b[16]) ;   // mult.v(2151)
    fa fa_17 (.a(wand_114), .b(wand_145), .cin(wand_176), .s(wfa_s_17), 
       .cout(wfa_cout_17));   // mult.v(2152)
    and (wand_207, a[6], b[15]) ;   // mult.v(2153)
    and (wand_238, a[7], b[14]) ;   // mult.v(2154)
    ha ha_7 (.a(wand_207), .b(wand_238), .s(wha_s_7), .c(wha_c_7));   // mult.v(2155)
    and (wand_22, a[0], b[22]) ;   // mult.v(2156)
    and (wand_53, a[1], b[21]) ;   // mult.v(2157)
    and (wand_84, a[2], b[20]) ;   // mult.v(2158)
    fa fa_18 (.a(wand_22), .b(wand_53), .cin(wand_84), .s(wfa_s_18), 
       .cout(wfa_cout_18));   // mult.v(2159)
    and (wand_115, a[3], b[19]) ;   // mult.v(2160)
    and (wand_146, a[4], b[18]) ;   // mult.v(2161)
    and (wand_177, a[5], b[17]) ;   // mult.v(2162)
    fa fa_19 (.a(wand_115), .b(wand_146), .cin(wand_177), .s(wfa_s_19), 
       .cout(wfa_cout_19));   // mult.v(2163)
    and (wand_208, a[6], b[16]) ;   // mult.v(2164)
    and (wand_239, a[7], b[15]) ;   // mult.v(2165)
    and (wand_270, a[8], b[14]) ;   // mult.v(2166)
    fa fa_20 (.a(wand_208), .b(wand_239), .cin(wand_270), .s(wfa_s_20), 
       .cout(wfa_cout_20));   // mult.v(2167)
    and (wand_301, a[9], b[13]) ;   // mult.v(2168)
    and (wand_332, a[10], b[12]) ;   // mult.v(2169)
    ha ha_8 (.a(wand_301), .b(wand_332), .s(wha_s_8), .c(wha_c_8));   // mult.v(2170)
    and (wand_23, a[0], b[23]) ;   // mult.v(2171)
    and (wand_54, a[1], b[22]) ;   // mult.v(2172)
    and (wand_85, a[2], b[21]) ;   // mult.v(2173)
    fa fa_21 (.a(wand_23), .b(wand_54), .cin(wand_85), .s(wfa_s_21), 
       .cout(wfa_cout_21));   // mult.v(2174)
    and (wand_116, a[3], b[20]) ;   // mult.v(2175)
    and (wand_147, a[4], b[19]) ;   // mult.v(2176)
    and (wand_178, a[5], b[18]) ;   // mult.v(2177)
    fa fa_22 (.a(wand_116), .b(wand_147), .cin(wand_178), .s(wfa_s_22), 
       .cout(wfa_cout_22));   // mult.v(2178)
    and (wand_209, a[6], b[17]) ;   // mult.v(2179)
    and (wand_240, a[7], b[16]) ;   // mult.v(2180)
    and (wand_271, a[8], b[15]) ;   // mult.v(2181)
    fa fa_23 (.a(wand_209), .b(wand_240), .cin(wand_271), .s(wfa_s_23), 
       .cout(wfa_cout_23));   // mult.v(2182)
    and (wand_302, a[9], b[14]) ;   // mult.v(2183)
    and (wand_333, a[10], b[13]) ;   // mult.v(2184)
    and (wand_364, a[11], b[12]) ;   // mult.v(2185)
    fa fa_24 (.a(wand_302), .b(wand_333), .cin(wand_364), .s(wfa_s_24), 
       .cout(wfa_cout_24));   // mult.v(2186)
    and (wand_395, a[12], b[11]) ;   // mult.v(2187)
    and (wand_426, a[13], b[10]) ;   // mult.v(2188)
    ha ha_9 (.a(wand_395), .b(wand_426), .s(wha_s_9), .c(wha_c_9));   // mult.v(2189)
    and (wand_24, a[0], b[24]) ;   // mult.v(2190)
    and (wand_55, a[1], b[23]) ;   // mult.v(2191)
    and (wand_86, a[2], b[22]) ;   // mult.v(2192)
    fa fa_25 (.a(wand_24), .b(wand_55), .cin(wand_86), .s(wfa_s_25), 
       .cout(wfa_cout_25));   // mult.v(2193)
    and (wand_117, a[3], b[21]) ;   // mult.v(2194)
    and (wand_148, a[4], b[20]) ;   // mult.v(2195)
    and (wand_179, a[5], b[19]) ;   // mult.v(2196)
    fa fa_26 (.a(wand_117), .b(wand_148), .cin(wand_179), .s(wfa_s_26), 
       .cout(wfa_cout_26));   // mult.v(2197)
    and (wand_210, a[6], b[18]) ;   // mult.v(2198)
    and (wand_241, a[7], b[17]) ;   // mult.v(2199)
    and (wand_272, a[8], b[16]) ;   // mult.v(2200)
    fa fa_27 (.a(wand_210), .b(wand_241), .cin(wand_272), .s(wfa_s_27), 
       .cout(wfa_cout_27));   // mult.v(2201)
    and (wand_303, a[9], b[15]) ;   // mult.v(2202)
    and (wand_334, a[10], b[14]) ;   // mult.v(2203)
    and (wand_365, a[11], b[13]) ;   // mult.v(2204)
    fa fa_28 (.a(wand_303), .b(wand_334), .cin(wand_365), .s(wfa_s_28), 
       .cout(wfa_cout_28));   // mult.v(2205)
    and (wand_396, a[12], b[12]) ;   // mult.v(2206)
    and (wand_427, a[13], b[11]) ;   // mult.v(2207)
    and (wand_458, a[14], b[10]) ;   // mult.v(2208)
    fa fa_29 (.a(wand_396), .b(wand_427), .cin(wand_458), .s(wfa_s_29), 
       .cout(wfa_cout_29));   // mult.v(2209)
    and (wand_489, a[15], b[9]) ;   // mult.v(2210)
    and (wand_520, a[16], b[8]) ;   // mult.v(2211)
    ha ha_10 (.a(wand_489), .b(wand_520), .s(wha_s_10), .c(wha_c_10));   // mult.v(2212)
    and (wand_25, a[0], b[25]) ;   // mult.v(2213)
    and (wand_56, a[1], b[24]) ;   // mult.v(2214)
    and (wand_87, a[2], b[23]) ;   // mult.v(2215)
    fa fa_30 (.a(wand_25), .b(wand_56), .cin(wand_87), .s(wfa_s_30), 
       .cout(wfa_cout_30));   // mult.v(2216)
    and (wand_118, a[3], b[22]) ;   // mult.v(2217)
    and (wand_149, a[4], b[21]) ;   // mult.v(2218)
    and (wand_180, a[5], b[20]) ;   // mult.v(2219)
    fa fa_31 (.a(wand_118), .b(wand_149), .cin(wand_180), .s(wfa_s_31), 
       .cout(wfa_cout_31));   // mult.v(2220)
    and (wand_211, a[6], b[19]) ;   // mult.v(2221)
    and (wand_242, a[7], b[18]) ;   // mult.v(2222)
    and (wand_273, a[8], b[17]) ;   // mult.v(2223)
    fa fa_32 (.a(wand_211), .b(wand_242), .cin(wand_273), .s(wfa_s_32), 
       .cout(wfa_cout_32));   // mult.v(2224)
    and (wand_304, a[9], b[16]) ;   // mult.v(2225)
    and (wand_335, a[10], b[15]) ;   // mult.v(2226)
    and (wand_366, a[11], b[14]) ;   // mult.v(2227)
    fa fa_33 (.a(wand_304), .b(wand_335), .cin(wand_366), .s(wfa_s_33), 
       .cout(wfa_cout_33));   // mult.v(2228)
    and (wand_397, a[12], b[13]) ;   // mult.v(2229)
    and (wand_428, a[13], b[12]) ;   // mult.v(2230)
    and (wand_459, a[14], b[11]) ;   // mult.v(2231)
    fa fa_34 (.a(wand_397), .b(wand_428), .cin(wand_459), .s(wfa_s_34), 
       .cout(wfa_cout_34));   // mult.v(2232)
    and (wand_490, a[15], b[10]) ;   // mult.v(2233)
    and (wand_521, a[16], b[9]) ;   // mult.v(2234)
    and (wand_552, a[17], b[8]) ;   // mult.v(2235)
    fa fa_35 (.a(wand_490), .b(wand_521), .cin(wand_552), .s(wfa_s_35), 
       .cout(wfa_cout_35));   // mult.v(2236)
    and (wand_583, a[18], b[7]) ;   // mult.v(2237)
    and (wand_614, a[19], b[6]) ;   // mult.v(2238)
    ha ha_11 (.a(wand_583), .b(wand_614), .s(wha_s_11), .c(wha_c_11));   // mult.v(2239)
    and (wand_26, a[0], b[26]) ;   // mult.v(2240)
    and (wand_57, a[1], b[25]) ;   // mult.v(2241)
    and (wand_88, a[2], b[24]) ;   // mult.v(2242)
    fa fa_36 (.a(wand_26), .b(wand_57), .cin(wand_88), .s(wfa_s_36), 
       .cout(wfa_cout_36));   // mult.v(2243)
    and (wand_119, a[3], b[23]) ;   // mult.v(2244)
    and (wand_150, a[4], b[22]) ;   // mult.v(2245)
    and (wand_181, a[5], b[21]) ;   // mult.v(2246)
    fa fa_37 (.a(wand_119), .b(wand_150), .cin(wand_181), .s(wfa_s_37), 
       .cout(wfa_cout_37));   // mult.v(2247)
    and (wand_212, a[6], b[20]) ;   // mult.v(2248)
    and (wand_243, a[7], b[19]) ;   // mult.v(2249)
    and (wand_274, a[8], b[18]) ;   // mult.v(2250)
    fa fa_38 (.a(wand_212), .b(wand_243), .cin(wand_274), .s(wfa_s_38), 
       .cout(wfa_cout_38));   // mult.v(2251)
    and (wand_305, a[9], b[17]) ;   // mult.v(2252)
    and (wand_336, a[10], b[16]) ;   // mult.v(2253)
    and (wand_367, a[11], b[15]) ;   // mult.v(2254)
    fa fa_39 (.a(wand_305), .b(wand_336), .cin(wand_367), .s(wfa_s_39), 
       .cout(wfa_cout_39));   // mult.v(2255)
    and (wand_398, a[12], b[14]) ;   // mult.v(2256)
    and (wand_429, a[13], b[13]) ;   // mult.v(2257)
    and (wand_460, a[14], b[12]) ;   // mult.v(2258)
    fa fa_40 (.a(wand_398), .b(wand_429), .cin(wand_460), .s(wfa_s_40), 
       .cout(wfa_cout_40));   // mult.v(2259)
    and (wand_491, a[15], b[11]) ;   // mult.v(2260)
    and (wand_522, a[16], b[10]) ;   // mult.v(2261)
    and (wand_553, a[17], b[9]) ;   // mult.v(2262)
    fa fa_41 (.a(wand_491), .b(wand_522), .cin(wand_553), .s(wfa_s_41), 
       .cout(wfa_cout_41));   // mult.v(2263)
    and (wand_584, a[18], b[8]) ;   // mult.v(2264)
    and (wand_615, a[19], b[7]) ;   // mult.v(2265)
    and (wand_646, a[20], b[6]) ;   // mult.v(2266)
    fa fa_42 (.a(wand_584), .b(wand_615), .cin(wand_646), .s(wfa_s_42), 
       .cout(wfa_cout_42));   // mult.v(2267)
    and (wand_677, a[21], b[5]) ;   // mult.v(2268)
    and (wand_708, a[22], b[4]) ;   // mult.v(2269)
    ha ha_12 (.a(wand_677), .b(wand_708), .s(wha_s_12), .c(wha_c_12));   // mult.v(2270)
    and (wand_27, a[0], b[27]) ;   // mult.v(2271)
    and (wand_58, a[1], b[26]) ;   // mult.v(2272)
    and (wand_89, a[2], b[25]) ;   // mult.v(2273)
    fa fa_43 (.a(wand_27), .b(wand_58), .cin(wand_89), .s(wfa_s_43), 
       .cout(wfa_cout_43));   // mult.v(2274)
    and (wand_120, a[3], b[24]) ;   // mult.v(2275)
    and (wand_151, a[4], b[23]) ;   // mult.v(2276)
    and (wand_182, a[5], b[22]) ;   // mult.v(2277)
    fa fa_44 (.a(wand_120), .b(wand_151), .cin(wand_182), .s(wfa_s_44), 
       .cout(wfa_cout_44));   // mult.v(2278)
    and (wand_213, a[6], b[21]) ;   // mult.v(2279)
    and (wand_244, a[7], b[20]) ;   // mult.v(2280)
    and (wand_275, a[8], b[19]) ;   // mult.v(2281)
    fa fa_45 (.a(wand_213), .b(wand_244), .cin(wand_275), .s(wfa_s_45), 
       .cout(wfa_cout_45));   // mult.v(2282)
    and (wand_306, a[9], b[18]) ;   // mult.v(2283)
    and (wand_337, a[10], b[17]) ;   // mult.v(2284)
    and (wand_368, a[11], b[16]) ;   // mult.v(2285)
    fa fa_46 (.a(wand_306), .b(wand_337), .cin(wand_368), .s(wfa_s_46), 
       .cout(wfa_cout_46));   // mult.v(2286)
    and (wand_399, a[12], b[15]) ;   // mult.v(2287)
    and (wand_430, a[13], b[14]) ;   // mult.v(2288)
    and (wand_461, a[14], b[13]) ;   // mult.v(2289)
    fa fa_47 (.a(wand_399), .b(wand_430), .cin(wand_461), .s(wfa_s_47), 
       .cout(wfa_cout_47));   // mult.v(2290)
    and (wand_492, a[15], b[12]) ;   // mult.v(2291)
    and (wand_523, a[16], b[11]) ;   // mult.v(2292)
    and (wand_554, a[17], b[10]) ;   // mult.v(2293)
    fa fa_48 (.a(wand_492), .b(wand_523), .cin(wand_554), .s(wfa_s_48), 
       .cout(wfa_cout_48));   // mult.v(2294)
    and (wand_585, a[18], b[9]) ;   // mult.v(2295)
    and (wand_616, a[19], b[8]) ;   // mult.v(2296)
    and (wand_647, a[20], b[7]) ;   // mult.v(2297)
    fa fa_49 (.a(wand_585), .b(wand_616), .cin(wand_647), .s(wfa_s_49), 
       .cout(wfa_cout_49));   // mult.v(2298)
    and (wand_678, a[21], b[6]) ;   // mult.v(2299)
    and (wand_709, a[22], b[5]) ;   // mult.v(2300)
    and (wand_740, a[23], b[4]) ;   // mult.v(2301)
    fa fa_50 (.a(wand_678), .b(wand_709), .cin(wand_740), .s(wfa_s_50), 
       .cout(wfa_cout_50));   // mult.v(2302)
    and (wand_771, a[24], b[3]) ;   // mult.v(2303)
    and (wand_802, a[25], b[2]) ;   // mult.v(2304)
    ha ha_13 (.a(wand_771), .b(wand_802), .s(wha_s_13), .c(wha_c_13));   // mult.v(2305)
    and (wand_90, a[2], b[26]) ;   // mult.v(2306)
    and (wand_121, a[3], b[25]) ;   // mult.v(2307)
    and (wand_152, a[4], b[24]) ;   // mult.v(2308)
    fa fa_51 (.a(wand_90), .b(wand_121), .cin(wand_152), .s(wfa_s_51), 
       .cout(wfa_cout_51));   // mult.v(2309)
    and (wand_183, a[5], b[23]) ;   // mult.v(2310)
    and (wand_214, a[6], b[22]) ;   // mult.v(2311)
    and (wand_245, a[7], b[21]) ;   // mult.v(2312)
    fa fa_52 (.a(wand_183), .b(wand_214), .cin(wand_245), .s(wfa_s_52), 
       .cout(wfa_cout_52));   // mult.v(2313)
    and (wand_276, a[8], b[20]) ;   // mult.v(2314)
    and (wand_307, a[9], b[19]) ;   // mult.v(2315)
    and (wand_338, a[10], b[18]) ;   // mult.v(2316)
    fa fa_53 (.a(wand_276), .b(wand_307), .cin(wand_338), .s(wfa_s_53), 
       .cout(wfa_cout_53));   // mult.v(2317)
    and (wand_369, a[11], b[17]) ;   // mult.v(2318)
    and (wand_400, a[12], b[16]) ;   // mult.v(2319)
    and (wand_431, a[13], b[15]) ;   // mult.v(2320)
    fa fa_54 (.a(wand_369), .b(wand_400), .cin(wand_431), .s(wfa_s_54), 
       .cout(wfa_cout_54));   // mult.v(2321)
    and (wand_462, a[14], b[14]) ;   // mult.v(2322)
    and (wand_493, a[15], b[13]) ;   // mult.v(2323)
    and (wand_524, a[16], b[12]) ;   // mult.v(2324)
    fa fa_55 (.a(wand_462), .b(wand_493), .cin(wand_524), .s(wfa_s_55), 
       .cout(wfa_cout_55));   // mult.v(2325)
    and (wand_555, a[17], b[11]) ;   // mult.v(2326)
    and (wand_586, a[18], b[10]) ;   // mult.v(2327)
    and (wand_617, a[19], b[9]) ;   // mult.v(2328)
    fa fa_56 (.a(wand_555), .b(wand_586), .cin(wand_617), .s(wfa_s_56), 
       .cout(wfa_cout_56));   // mult.v(2329)
    and (wand_648, a[20], b[8]) ;   // mult.v(2330)
    and (wand_679, a[21], b[7]) ;   // mult.v(2331)
    and (wand_710, a[22], b[6]) ;   // mult.v(2332)
    fa fa_57 (.a(wand_648), .b(wand_679), .cin(wand_710), .s(wfa_s_57), 
       .cout(wfa_cout_57));   // mult.v(2333)
    and (wand_741, a[23], b[5]) ;   // mult.v(2334)
    and (wand_772, a[24], b[4]) ;   // mult.v(2335)
    and (wand_803, a[25], b[3]) ;   // mult.v(2336)
    fa fa_58 (.a(wand_741), .b(wand_772), .cin(wand_803), .s(wfa_s_58), 
       .cout(wfa_cout_58));   // mult.v(2337)
    and (wand_834, a[26], b[2]) ;   // mult.v(2338)
    and (wand_865, a[27], b[1]) ;   // mult.v(2339)
    and (wand_896, a[28], b[0]) ;   // mult.v(2340)
    fa fa_59 (.a(wand_834), .b(wand_865), .cin(wand_896), .s(wfa_s_59), 
       .cout(wfa_cout_59));   // mult.v(2341)
    and (wand_184, a[5], b[24]) ;   // mult.v(2342)
    and (wand_215, a[6], b[23]) ;   // mult.v(2343)
    and (wand_246, a[7], b[22]) ;   // mult.v(2344)
    fa fa_60 (.a(wand_184), .b(wand_215), .cin(wand_246), .s(wfa_s_60), 
       .cout(wfa_cout_60));   // mult.v(2345)
    and (wand_277, a[8], b[21]) ;   // mult.v(2346)
    and (wand_308, a[9], b[20]) ;   // mult.v(2347)
    and (wand_339, a[10], b[19]) ;   // mult.v(2348)
    fa fa_61 (.a(wand_277), .b(wand_308), .cin(wand_339), .s(wfa_s_61), 
       .cout(wfa_cout_61));   // mult.v(2349)
    and (wand_370, a[11], b[18]) ;   // mult.v(2350)
    and (wand_401, a[12], b[17]) ;   // mult.v(2351)
    and (wand_432, a[13], b[16]) ;   // mult.v(2352)
    fa fa_62 (.a(wand_370), .b(wand_401), .cin(wand_432), .s(wfa_s_62), 
       .cout(wfa_cout_62));   // mult.v(2353)
    and (wand_463, a[14], b[15]) ;   // mult.v(2354)
    and (wand_494, a[15], b[14]) ;   // mult.v(2355)
    and (wand_525, a[16], b[13]) ;   // mult.v(2356)
    fa fa_63 (.a(wand_463), .b(wand_494), .cin(wand_525), .s(wfa_s_63), 
       .cout(wfa_cout_63));   // mult.v(2357)
    and (wand_556, a[17], b[12]) ;   // mult.v(2358)
    and (wand_587, a[18], b[11]) ;   // mult.v(2359)
    and (wand_618, a[19], b[10]) ;   // mult.v(2360)
    fa fa_64 (.a(wand_556), .b(wand_587), .cin(wand_618), .s(wfa_s_64), 
       .cout(wfa_cout_64));   // mult.v(2361)
    and (wand_649, a[20], b[9]) ;   // mult.v(2362)
    and (wand_680, a[21], b[8]) ;   // mult.v(2363)
    and (wand_711, a[22], b[7]) ;   // mult.v(2364)
    fa fa_65 (.a(wand_649), .b(wand_680), .cin(wand_711), .s(wfa_s_65), 
       .cout(wfa_cout_65));   // mult.v(2365)
    and (wand_742, a[23], b[6]) ;   // mult.v(2366)
    and (wand_773, a[24], b[5]) ;   // mult.v(2367)
    and (wand_804, a[25], b[4]) ;   // mult.v(2368)
    fa fa_66 (.a(wand_742), .b(wand_773), .cin(wand_804), .s(wfa_s_66), 
       .cout(wfa_cout_66));   // mult.v(2369)
    and (wand_835, a[26], b[3]) ;   // mult.v(2370)
    and (wand_866, a[27], b[2]) ;   // mult.v(2371)
    and (wand_897, a[28], b[1]) ;   // mult.v(2372)
    fa fa_67 (.a(wand_835), .b(wand_866), .cin(wand_897), .s(wfa_s_67), 
       .cout(wfa_cout_67));   // mult.v(2373)
    and (wand_928, a[29], b[0]) ;   // mult.v(2374)
    fa fa_68 (.a(wand_928), .b(wha_c_0), .cin(wfa_s_0), .s(wfa_s_68), 
       .cout(wfa_cout_68));   // mult.v(2375)
    and (wand_278, a[8], b[22]) ;   // mult.v(2376)
    and (wand_309, a[9], b[21]) ;   // mult.v(2377)
    and (wand_340, a[10], b[20]) ;   // mult.v(2378)
    fa fa_69 (.a(wand_278), .b(wand_309), .cin(wand_340), .s(wfa_s_69), 
       .cout(wfa_cout_69));   // mult.v(2379)
    and (wand_371, a[11], b[19]) ;   // mult.v(2380)
    and (wand_402, a[12], b[18]) ;   // mult.v(2381)
    and (wand_433, a[13], b[17]) ;   // mult.v(2382)
    fa fa_70 (.a(wand_371), .b(wand_402), .cin(wand_433), .s(wfa_s_70), 
       .cout(wfa_cout_70));   // mult.v(2383)
    and (wand_464, a[14], b[16]) ;   // mult.v(2384)
    and (wand_495, a[15], b[15]) ;   // mult.v(2385)
    and (wand_526, a[16], b[14]) ;   // mult.v(2386)
    fa fa_71 (.a(wand_464), .b(wand_495), .cin(wand_526), .s(wfa_s_71), 
       .cout(wfa_cout_71));   // mult.v(2387)
    and (wand_557, a[17], b[13]) ;   // mult.v(2388)
    and (wand_588, a[18], b[12]) ;   // mult.v(2389)
    and (wand_619, a[19], b[11]) ;   // mult.v(2390)
    fa fa_72 (.a(wand_557), .b(wand_588), .cin(wand_619), .s(wfa_s_72), 
       .cout(wfa_cout_72));   // mult.v(2391)
    and (wand_650, a[20], b[10]) ;   // mult.v(2392)
    and (wand_681, a[21], b[9]) ;   // mult.v(2393)
    and (wand_712, a[22], b[8]) ;   // mult.v(2394)
    fa fa_73 (.a(wand_650), .b(wand_681), .cin(wand_712), .s(wfa_s_73), 
       .cout(wfa_cout_73));   // mult.v(2395)
    and (wand_743, a[23], b[7]) ;   // mult.v(2396)
    and (wand_774, a[24], b[6]) ;   // mult.v(2397)
    and (wand_805, a[25], b[5]) ;   // mult.v(2398)
    fa fa_74 (.a(wand_743), .b(wand_774), .cin(wand_805), .s(wfa_s_74), 
       .cout(wfa_cout_74));   // mult.v(2399)
    and (wand_836, a[26], b[4]) ;   // mult.v(2400)
    and (wand_867, a[27], b[3]) ;   // mult.v(2401)
    and (wand_898, a[28], b[2]) ;   // mult.v(2402)
    fa fa_75 (.a(wand_836), .b(wand_867), .cin(wand_898), .s(wfa_s_75), 
       .cout(wfa_cout_75));   // mult.v(2403)
    and (wand_929, a[29], b[1]) ;   // mult.v(2404)
    and (wand_960, a[30], b[0]) ;   // mult.v(2405)
    fa fa_76 (.a(wand_929), .b(wand_960), .cin(wfa_cout_0), .s(wfa_s_76), 
       .cout(wfa_cout_76));   // mult.v(2406)
    fa fa_77 (.a(wha_c_1), .b(wfa_s_1), .cin(wfa_s_2), .s(wfa_s_77), 
       .cout(wfa_cout_77));   // mult.v(2407)
    and (wand_372, a[11], b[20]) ;   // mult.v(2408)
    and (wand_403, a[12], b[19]) ;   // mult.v(2409)
    and (wand_434, a[13], b[18]) ;   // mult.v(2410)
    fa fa_78 (.a(wand_372), .b(wand_403), .cin(wand_434), .s(wfa_s_78), 
       .cout(wfa_cout_78));   // mult.v(2411)
    and (wand_465, a[14], b[17]) ;   // mult.v(2412)
    and (wand_496, a[15], b[16]) ;   // mult.v(2413)
    and (wand_527, a[16], b[15]) ;   // mult.v(2414)
    fa fa_79 (.a(wand_465), .b(wand_496), .cin(wand_527), .s(wfa_s_79), 
       .cout(wfa_cout_79));   // mult.v(2415)
    and (wand_558, a[17], b[14]) ;   // mult.v(2416)
    and (wand_589, a[18], b[13]) ;   // mult.v(2417)
    and (wand_620, a[19], b[12]) ;   // mult.v(2418)
    fa fa_80 (.a(wand_558), .b(wand_589), .cin(wand_620), .s(wfa_s_80), 
       .cout(wfa_cout_80));   // mult.v(2419)
    and (wand_651, a[20], b[11]) ;   // mult.v(2420)
    and (wand_682, a[21], b[10]) ;   // mult.v(2421)
    and (wand_713, a[22], b[9]) ;   // mult.v(2422)
    fa fa_81 (.a(wand_651), .b(wand_682), .cin(wand_713), .s(wfa_s_81), 
       .cout(wfa_cout_81));   // mult.v(2423)
    and (wand_744, a[23], b[8]) ;   // mult.v(2424)
    and (wand_775, a[24], b[7]) ;   // mult.v(2425)
    and (wand_806, a[25], b[6]) ;   // mult.v(2426)
    fa fa_82 (.a(wand_744), .b(wand_775), .cin(wand_806), .s(wfa_s_82), 
       .cout(wfa_cout_82));   // mult.v(2427)
    and (wand_837, a[26], b[5]) ;   // mult.v(2428)
    and (wand_868, a[27], b[4]) ;   // mult.v(2429)
    and (wand_899, a[28], b[3]) ;   // mult.v(2430)
    fa fa_83 (.a(wand_837), .b(wand_868), .cin(wand_899), .s(wfa_s_83), 
       .cout(wfa_cout_83));   // mult.v(2431)
    and (wand_930, a[29], b[2]) ;   // mult.v(2432)
    and (wand_961, a[30], b[1]) ;   // mult.v(2433)
    and (wand_992, a[31], b[0]) ;   // mult.v(2434)
    fa fa_84 (.a(wand_930), .b(wand_961), .cin(wand_992), .s(wfa_s_84), 
       .cout(wfa_cout_84));   // mult.v(2435)
    fa fa_85 (.a(wfa_cout_1), .b(wfa_cout_2), .cin(wha_c_2), .s(wfa_s_85), 
       .cout(wfa_cout_85));   // mult.v(2436)
    fa fa_86 (.a(wfa_s_3), .b(wfa_s_4), .cin(wfa_s_5), .s(wfa_s_86), 
       .cout(wfa_cout_86));   // mult.v(2437)
    and (wand_404, a[12], b[20]) ;   // mult.v(2438)
    and (wand_435, a[13], b[19]) ;   // mult.v(2439)
    and (wand_466, a[14], b[18]) ;   // mult.v(2440)
    fa fa_87 (.a(wand_404), .b(wand_435), .cin(wand_466), .s(wfa_s_87), 
       .cout(wfa_cout_87));   // mult.v(2441)
    and (wand_497, a[15], b[17]) ;   // mult.v(2442)
    and (wand_528, a[16], b[16]) ;   // mult.v(2443)
    and (wand_559, a[17], b[15]) ;   // mult.v(2444)
    fa fa_88 (.a(wand_497), .b(wand_528), .cin(wand_559), .s(wfa_s_88), 
       .cout(wfa_cout_88));   // mult.v(2445)
    and (wand_590, a[18], b[14]) ;   // mult.v(2446)
    and (wand_621, a[19], b[13]) ;   // mult.v(2447)
    and (wand_652, a[20], b[12]) ;   // mult.v(2448)
    fa fa_89 (.a(wand_590), .b(wand_621), .cin(wand_652), .s(wfa_s_89), 
       .cout(wfa_cout_89));   // mult.v(2449)
    and (wand_683, a[21], b[11]) ;   // mult.v(2450)
    and (wand_714, a[22], b[10]) ;   // mult.v(2451)
    and (wand_745, a[23], b[9]) ;   // mult.v(2452)
    fa fa_90 (.a(wand_683), .b(wand_714), .cin(wand_745), .s(wfa_s_90), 
       .cout(wfa_cout_90));   // mult.v(2453)
    and (wand_776, a[24], b[8]) ;   // mult.v(2454)
    and (wand_807, a[25], b[7]) ;   // mult.v(2455)
    and (wand_838, a[26], b[6]) ;   // mult.v(2456)
    fa fa_91 (.a(wand_776), .b(wand_807), .cin(wand_838), .s(wfa_s_91), 
       .cout(wfa_cout_91));   // mult.v(2457)
    and (wand_869, a[27], b[5]) ;   // mult.v(2458)
    and (wand_900, a[28], b[4]) ;   // mult.v(2459)
    and (wand_931, a[29], b[3]) ;   // mult.v(2460)
    fa fa_92 (.a(wand_869), .b(wand_900), .cin(wand_931), .s(wfa_s_92), 
       .cout(wfa_cout_92));   // mult.v(2461)
    and (wand_962, a[30], b[2]) ;   // mult.v(2462)
    and (wand_993, a[31], b[1]) ;   // mult.v(2463)
    fa fa_93 (.a(wand_962), .b(wand_993), .cin(wfa_cout_3), .s(wfa_s_93), 
       .cout(wfa_cout_93));   // mult.v(2464)
    fa fa_94 (.a(wfa_cout_4), .b(wfa_cout_5), .cin(wha_c_3), .s(wfa_s_94), 
       .cout(wfa_cout_94));   // mult.v(2465)
    fa fa_95 (.a(wfa_s_6), .b(wfa_s_7), .cin(wfa_s_8), .s(wfa_s_95), 
       .cout(wfa_cout_95));   // mult.v(2466)
    and (wand_374, a[11], b[22]) ;   // mult.v(2467)
    and (wand_405, a[12], b[21]) ;   // mult.v(2468)
    and (wand_436, a[13], b[20]) ;   // mult.v(2469)
    fa fa_96 (.a(wand_374), .b(wand_405), .cin(wand_436), .s(wfa_s_96), 
       .cout(wfa_cout_96));   // mult.v(2470)
    and (wand_467, a[14], b[19]) ;   // mult.v(2471)
    and (wand_498, a[15], b[18]) ;   // mult.v(2472)
    and (wand_529, a[16], b[17]) ;   // mult.v(2473)
    fa fa_97 (.a(wand_467), .b(wand_498), .cin(wand_529), .s(wfa_s_97), 
       .cout(wfa_cout_97));   // mult.v(2474)
    and (wand_560, a[17], b[16]) ;   // mult.v(2475)
    and (wand_591, a[18], b[15]) ;   // mult.v(2476)
    and (wand_622, a[19], b[14]) ;   // mult.v(2477)
    fa fa_98 (.a(wand_560), .b(wand_591), .cin(wand_622), .s(wfa_s_98), 
       .cout(wfa_cout_98));   // mult.v(2478)
    and (wand_653, a[20], b[13]) ;   // mult.v(2479)
    and (wand_684, a[21], b[12]) ;   // mult.v(2480)
    and (wand_715, a[22], b[11]) ;   // mult.v(2481)
    fa fa_99 (.a(wand_653), .b(wand_684), .cin(wand_715), .s(wfa_s_99), 
       .cout(wfa_cout_99));   // mult.v(2482)
    and (wand_746, a[23], b[10]) ;   // mult.v(2483)
    and (wand_777, a[24], b[9]) ;   // mult.v(2484)
    and (wand_808, a[25], b[8]) ;   // mult.v(2485)
    fa fa_100 (.a(wand_746), .b(wand_777), .cin(wand_808), .s(wfa_s_100), 
       .cout(wfa_cout_100));   // mult.v(2486)
    and (wand_839, a[26], b[7]) ;   // mult.v(2487)
    and (wand_870, a[27], b[6]) ;   // mult.v(2488)
    and (wand_901, a[28], b[5]) ;   // mult.v(2489)
    fa fa_101 (.a(wand_839), .b(wand_870), .cin(wand_901), .s(wfa_s_101), 
       .cout(wfa_cout_101));   // mult.v(2490)
    and (wand_932, a[29], b[4]) ;   // mult.v(2491)
    and (wand_963, a[30], b[3]) ;   // mult.v(2492)
    and (wand_994, a[31], b[2]) ;   // mult.v(2493)
    fa fa_102 (.a(wand_932), .b(wand_963), .cin(wand_994), .s(wfa_s_102), 
       .cout(wfa_cout_102));   // mult.v(2494)
    fa fa_103 (.a(wfa_cout_6), .b(wfa_cout_7), .cin(wfa_cout_8), .s(wfa_s_103), 
       .cout(wfa_cout_103));   // mult.v(2495)
    fa fa_104 (.a(wha_c_4), .b(wfa_s_9), .cin(wfa_s_10), .s(wfa_s_104), 
       .cout(wfa_cout_104));   // mult.v(2496)
    and (wand_313, a[9], b[25]) ;   // mult.v(2497)
    and (wand_344, a[10], b[24]) ;   // mult.v(2498)
    and (wand_375, a[11], b[23]) ;   // mult.v(2499)
    fa fa_105 (.a(wand_313), .b(wand_344), .cin(wand_375), .s(wfa_s_105), 
       .cout(wfa_cout_105));   // mult.v(2500)
    and (wand_406, a[12], b[22]) ;   // mult.v(2501)
    and (wand_437, a[13], b[21]) ;   // mult.v(2502)
    and (wand_468, a[14], b[20]) ;   // mult.v(2503)
    fa fa_106 (.a(wand_406), .b(wand_437), .cin(wand_468), .s(wfa_s_106), 
       .cout(wfa_cout_106));   // mult.v(2504)
    and (wand_499, a[15], b[19]) ;   // mult.v(2505)
    and (wand_530, a[16], b[18]) ;   // mult.v(2506)
    and (wand_561, a[17], b[17]) ;   // mult.v(2507)
    fa fa_107 (.a(wand_499), .b(wand_530), .cin(wand_561), .s(wfa_s_107), 
       .cout(wfa_cout_107));   // mult.v(2508)
    and (wand_592, a[18], b[16]) ;   // mult.v(2509)
    and (wand_623, a[19], b[15]) ;   // mult.v(2510)
    and (wand_654, a[20], b[14]) ;   // mult.v(2511)
    fa fa_108 (.a(wand_592), .b(wand_623), .cin(wand_654), .s(wfa_s_108), 
       .cout(wfa_cout_108));   // mult.v(2512)
    and (wand_685, a[21], b[13]) ;   // mult.v(2513)
    and (wand_716, a[22], b[12]) ;   // mult.v(2514)
    and (wand_747, a[23], b[11]) ;   // mult.v(2515)
    fa fa_109 (.a(wand_685), .b(wand_716), .cin(wand_747), .s(wfa_s_109), 
       .cout(wfa_cout_109));   // mult.v(2516)
    and (wand_778, a[24], b[10]) ;   // mult.v(2517)
    and (wand_809, a[25], b[9]) ;   // mult.v(2518)
    and (wand_840, a[26], b[8]) ;   // mult.v(2519)
    fa fa_110 (.a(wand_778), .b(wand_809), .cin(wand_840), .s(wfa_s_110), 
       .cout(wfa_cout_110));   // mult.v(2520)
    and (wand_871, a[27], b[7]) ;   // mult.v(2521)
    and (wand_902, a[28], b[6]) ;   // mult.v(2522)
    and (wand_933, a[29], b[5]) ;   // mult.v(2523)
    fa fa_111 (.a(wand_871), .b(wand_902), .cin(wand_933), .s(wfa_s_111), 
       .cout(wfa_cout_111));   // mult.v(2524)
    and (wand_964, a[30], b[4]) ;   // mult.v(2525)
    and (wand_995, a[31], b[3]) ;   // mult.v(2526)
    fa fa_112 (.a(wand_964), .b(wand_995), .cin(wfa_cout_9), .s(wfa_s_112), 
       .cout(wfa_cout_112));   // mult.v(2527)
    fa fa_113 (.a(wfa_cout_10), .b(wfa_cout_11), .cin(wfa_s_12), .s(wfa_s_113), 
       .cout(wfa_cout_113));   // mult.v(2528)
    and (wand_252, a[7], b[28]) ;   // mult.v(2529)
    and (wand_283, a[8], b[27]) ;   // mult.v(2530)
    and (wand_314, a[9], b[26]) ;   // mult.v(2531)
    fa fa_114 (.a(wand_252), .b(wand_283), .cin(wand_314), .s(wfa_s_114), 
       .cout(wfa_cout_114));   // mult.v(2532)
    and (wand_345, a[10], b[25]) ;   // mult.v(2533)
    and (wand_376, a[11], b[24]) ;   // mult.v(2534)
    and (wand_407, a[12], b[23]) ;   // mult.v(2535)
    fa fa_115 (.a(wand_345), .b(wand_376), .cin(wand_407), .s(wfa_s_115), 
       .cout(wfa_cout_115));   // mult.v(2536)
    and (wand_438, a[13], b[22]) ;   // mult.v(2537)
    and (wand_469, a[14], b[21]) ;   // mult.v(2538)
    and (wand_500, a[15], b[20]) ;   // mult.v(2539)
    fa fa_116 (.a(wand_438), .b(wand_469), .cin(wand_500), .s(wfa_s_116), 
       .cout(wfa_cout_116));   // mult.v(2540)
    and (wand_531, a[16], b[19]) ;   // mult.v(2541)
    and (wand_562, a[17], b[18]) ;   // mult.v(2542)
    and (wand_593, a[18], b[17]) ;   // mult.v(2543)
    fa fa_117 (.a(wand_531), .b(wand_562), .cin(wand_593), .s(wfa_s_117), 
       .cout(wfa_cout_117));   // mult.v(2544)
    and (wand_624, a[19], b[16]) ;   // mult.v(2545)
    and (wand_655, a[20], b[15]) ;   // mult.v(2546)
    and (wand_686, a[21], b[14]) ;   // mult.v(2547)
    fa fa_118 (.a(wand_624), .b(wand_655), .cin(wand_686), .s(wfa_s_118), 
       .cout(wfa_cout_118));   // mult.v(2548)
    and (wand_717, a[22], b[13]) ;   // mult.v(2549)
    and (wand_748, a[23], b[12]) ;   // mult.v(2550)
    and (wand_779, a[24], b[11]) ;   // mult.v(2551)
    fa fa_119 (.a(wand_717), .b(wand_748), .cin(wand_779), .s(wfa_s_119), 
       .cout(wfa_cout_119));   // mult.v(2552)
    and (wand_810, a[25], b[10]) ;   // mult.v(2553)
    and (wand_841, a[26], b[9]) ;   // mult.v(2554)
    and (wand_872, a[27], b[8]) ;   // mult.v(2555)
    fa fa_120 (.a(wand_810), .b(wand_841), .cin(wand_872), .s(wfa_s_120), 
       .cout(wfa_cout_120));   // mult.v(2556)
    and (wand_903, a[28], b[7]) ;   // mult.v(2557)
    and (wand_934, a[29], b[6]) ;   // mult.v(2558)
    and (wand_965, a[30], b[5]) ;   // mult.v(2559)
    fa fa_121 (.a(wand_903), .b(wand_934), .cin(wand_965), .s(wfa_s_121), 
       .cout(wfa_cout_121));   // mult.v(2560)
    and (wand_996, a[31], b[4]) ;   // mult.v(2561)
    fa fa_122 (.a(wand_996), .b(wfa_cout_12), .cin(wfa_cout_13), .s(wfa_s_122), 
       .cout(wfa_cout_122));   // mult.v(2562)
    and (wand_191, a[5], b[31]) ;   // mult.v(2563)
    and (wand_222, a[6], b[30]) ;   // mult.v(2564)
    and (wand_253, a[7], b[29]) ;   // mult.v(2565)
    fa fa_123 (.a(wand_191), .b(wand_222), .cin(wand_253), .s(wfa_s_123), 
       .cout(wfa_cout_123));   // mult.v(2566)
    and (wand_284, a[8], b[28]) ;   // mult.v(2567)
    and (wand_315, a[9], b[27]) ;   // mult.v(2568)
    and (wand_346, a[10], b[26]) ;   // mult.v(2569)
    fa fa_124 (.a(wand_284), .b(wand_315), .cin(wand_346), .s(wfa_s_124), 
       .cout(wfa_cout_124));   // mult.v(2570)
    and (wand_377, a[11], b[25]) ;   // mult.v(2571)
    and (wand_408, a[12], b[24]) ;   // mult.v(2572)
    and (wand_439, a[13], b[23]) ;   // mult.v(2573)
    fa fa_125 (.a(wand_377), .b(wand_408), .cin(wand_439), .s(wfa_s_125), 
       .cout(wfa_cout_125));   // mult.v(2574)
    and (wand_470, a[14], b[22]) ;   // mult.v(2575)
    and (wand_501, a[15], b[21]) ;   // mult.v(2576)
    and (wand_532, a[16], b[20]) ;   // mult.v(2577)
    fa fa_126 (.a(wand_470), .b(wand_501), .cin(wand_532), .s(wfa_s_126), 
       .cout(wfa_cout_126));   // mult.v(2578)
    and (wand_563, a[17], b[19]) ;   // mult.v(2579)
    and (wand_594, a[18], b[18]) ;   // mult.v(2580)
    and (wand_625, a[19], b[17]) ;   // mult.v(2581)
    fa fa_127 (.a(wand_563), .b(wand_594), .cin(wand_625), .s(wfa_s_127), 
       .cout(wfa_cout_127));   // mult.v(2582)
    and (wand_656, a[20], b[16]) ;   // mult.v(2583)
    and (wand_687, a[21], b[15]) ;   // mult.v(2584)
    and (wand_718, a[22], b[14]) ;   // mult.v(2585)
    fa fa_128 (.a(wand_656), .b(wand_687), .cin(wand_718), .s(wfa_s_128), 
       .cout(wfa_cout_128));   // mult.v(2586)
    and (wand_749, a[23], b[13]) ;   // mult.v(2587)
    and (wand_780, a[24], b[12]) ;   // mult.v(2588)
    and (wand_811, a[25], b[11]) ;   // mult.v(2589)
    fa fa_129 (.a(wand_749), .b(wand_780), .cin(wand_811), .s(wfa_s_129), 
       .cout(wfa_cout_129));   // mult.v(2590)
    and (wand_842, a[26], b[10]) ;   // mult.v(2591)
    and (wand_873, a[27], b[9]) ;   // mult.v(2592)
    and (wand_904, a[28], b[8]) ;   // mult.v(2593)
    fa fa_130 (.a(wand_842), .b(wand_873), .cin(wand_904), .s(wfa_s_130), 
       .cout(wfa_cout_130));   // mult.v(2594)
    and (wand_935, a[29], b[7]) ;   // mult.v(2595)
    and (wand_966, a[30], b[6]) ;   // mult.v(2596)
    and (wand_997, a[31], b[5]) ;   // mult.v(2597)
    fa fa_131 (.a(wand_935), .b(wand_966), .cin(wand_997), .s(wfa_s_131), 
       .cout(wfa_cout_131));   // mult.v(2598)
    and (wand_223, a[6], b[31]) ;   // mult.v(2599)
    and (wand_254, a[7], b[30]) ;   // mult.v(2600)
    and (wand_285, a[8], b[29]) ;   // mult.v(2601)
    fa fa_132 (.a(wand_223), .b(wand_254), .cin(wand_285), .s(wfa_s_132), 
       .cout(wfa_cout_132));   // mult.v(2602)
    and (wand_316, a[9], b[28]) ;   // mult.v(2603)
    and (wand_347, a[10], b[27]) ;   // mult.v(2604)
    and (wand_378, a[11], b[26]) ;   // mult.v(2605)
    fa fa_133 (.a(wand_316), .b(wand_347), .cin(wand_378), .s(wfa_s_133), 
       .cout(wfa_cout_133));   // mult.v(2606)
    and (wand_409, a[12], b[25]) ;   // mult.v(2607)
    and (wand_440, a[13], b[24]) ;   // mult.v(2608)
    and (wand_471, a[14], b[23]) ;   // mult.v(2609)
    fa fa_134 (.a(wand_409), .b(wand_440), .cin(wand_471), .s(wfa_s_134), 
       .cout(wfa_cout_134));   // mult.v(2610)
    and (wand_502, a[15], b[22]) ;   // mult.v(2611)
    and (wand_533, a[16], b[21]) ;   // mult.v(2612)
    and (wand_564, a[17], b[20]) ;   // mult.v(2613)
    fa fa_135 (.a(wand_502), .b(wand_533), .cin(wand_564), .s(wfa_s_135), 
       .cout(wfa_cout_135));   // mult.v(2614)
    and (wand_595, a[18], b[19]) ;   // mult.v(2615)
    and (wand_626, a[19], b[18]) ;   // mult.v(2616)
    and (wand_657, a[20], b[17]) ;   // mult.v(2617)
    fa fa_136 (.a(wand_595), .b(wand_626), .cin(wand_657), .s(wfa_s_136), 
       .cout(wfa_cout_136));   // mult.v(2618)
    and (wand_688, a[21], b[16]) ;   // mult.v(2619)
    and (wand_719, a[22], b[15]) ;   // mult.v(2620)
    and (wand_750, a[23], b[14]) ;   // mult.v(2621)
    fa fa_137 (.a(wand_688), .b(wand_719), .cin(wand_750), .s(wfa_s_137), 
       .cout(wfa_cout_137));   // mult.v(2622)
    and (wand_781, a[24], b[13]) ;   // mult.v(2623)
    and (wand_812, a[25], b[12]) ;   // mult.v(2624)
    and (wand_843, a[26], b[11]) ;   // mult.v(2625)
    fa fa_138 (.a(wand_781), .b(wand_812), .cin(wand_843), .s(wfa_s_138), 
       .cout(wfa_cout_138));   // mult.v(2626)
    and (wand_874, a[27], b[10]) ;   // mult.v(2627)
    and (wand_905, a[28], b[9]) ;   // mult.v(2628)
    and (wand_936, a[29], b[8]) ;   // mult.v(2629)
    fa fa_139 (.a(wand_874), .b(wand_905), .cin(wand_936), .s(wfa_s_139), 
       .cout(wfa_cout_139));   // mult.v(2630)
    and (wand_255, a[7], b[31]) ;   // mult.v(2631)
    and (wand_286, a[8], b[30]) ;   // mult.v(2632)
    and (wand_317, a[9], b[29]) ;   // mult.v(2633)
    fa fa_140 (.a(wand_255), .b(wand_286), .cin(wand_317), .s(wfa_s_140), 
       .cout(wfa_cout_140));   // mult.v(2634)
    and (wand_348, a[10], b[28]) ;   // mult.v(2635)
    and (wand_379, a[11], b[27]) ;   // mult.v(2636)
    and (wand_410, a[12], b[26]) ;   // mult.v(2637)
    fa fa_141 (.a(wand_348), .b(wand_379), .cin(wand_410), .s(wfa_s_141), 
       .cout(wfa_cout_141));   // mult.v(2638)
    and (wand_441, a[13], b[25]) ;   // mult.v(2639)
    and (wand_472, a[14], b[24]) ;   // mult.v(2640)
    and (wand_503, a[15], b[23]) ;   // mult.v(2641)
    fa fa_142 (.a(wand_441), .b(wand_472), .cin(wand_503), .s(wfa_s_142), 
       .cout(wfa_cout_142));   // mult.v(2642)
    and (wand_534, a[16], b[22]) ;   // mult.v(2643)
    and (wand_565, a[17], b[21]) ;   // mult.v(2644)
    and (wand_596, a[18], b[20]) ;   // mult.v(2645)
    fa fa_143 (.a(wand_534), .b(wand_565), .cin(wand_596), .s(wfa_s_143), 
       .cout(wfa_cout_143));   // mult.v(2646)
    and (wand_627, a[19], b[19]) ;   // mult.v(2647)
    and (wand_658, a[20], b[18]) ;   // mult.v(2648)
    and (wand_689, a[21], b[17]) ;   // mult.v(2649)
    fa fa_144 (.a(wand_627), .b(wand_658), .cin(wand_689), .s(wfa_s_144), 
       .cout(wfa_cout_144));   // mult.v(2650)
    and (wand_720, a[22], b[16]) ;   // mult.v(2651)
    and (wand_751, a[23], b[15]) ;   // mult.v(2652)
    and (wand_782, a[24], b[14]) ;   // mult.v(2653)
    fa fa_145 (.a(wand_720), .b(wand_751), .cin(wand_782), .s(wfa_s_145), 
       .cout(wfa_cout_145));   // mult.v(2654)
    and (wand_813, a[25], b[13]) ;   // mult.v(2655)
    and (wand_844, a[26], b[12]) ;   // mult.v(2656)
    and (wand_875, a[27], b[11]) ;   // mult.v(2657)
    fa fa_146 (.a(wand_813), .b(wand_844), .cin(wand_875), .s(wfa_s_146), 
       .cout(wfa_cout_146));   // mult.v(2658)
    and (wand_287, a[8], b[31]) ;   // mult.v(2659)
    and (wand_318, a[9], b[30]) ;   // mult.v(2660)
    and (wand_349, a[10], b[29]) ;   // mult.v(2661)
    fa fa_147 (.a(wand_287), .b(wand_318), .cin(wand_349), .s(wfa_s_147), 
       .cout(wfa_cout_147));   // mult.v(2662)
    and (wand_380, a[11], b[28]) ;   // mult.v(2663)
    and (wand_411, a[12], b[27]) ;   // mult.v(2664)
    and (wand_442, a[13], b[26]) ;   // mult.v(2665)
    fa fa_148 (.a(wand_380), .b(wand_411), .cin(wand_442), .s(wfa_s_148), 
       .cout(wfa_cout_148));   // mult.v(2666)
    and (wand_473, a[14], b[25]) ;   // mult.v(2667)
    and (wand_504, a[15], b[24]) ;   // mult.v(2668)
    and (wand_535, a[16], b[23]) ;   // mult.v(2669)
    fa fa_149 (.a(wand_473), .b(wand_504), .cin(wand_535), .s(wfa_s_149), 
       .cout(wfa_cout_149));   // mult.v(2670)
    and (wand_566, a[17], b[22]) ;   // mult.v(2671)
    and (wand_597, a[18], b[21]) ;   // mult.v(2672)
    and (wand_628, a[19], b[20]) ;   // mult.v(2673)
    fa fa_150 (.a(wand_566), .b(wand_597), .cin(wand_628), .s(wfa_s_150), 
       .cout(wfa_cout_150));   // mult.v(2674)
    and (wand_659, a[20], b[19]) ;   // mult.v(2675)
    and (wand_690, a[21], b[18]) ;   // mult.v(2676)
    and (wand_721, a[22], b[17]) ;   // mult.v(2677)
    fa fa_151 (.a(wand_659), .b(wand_690), .cin(wand_721), .s(wfa_s_151), 
       .cout(wfa_cout_151));   // mult.v(2678)
    and (wand_752, a[23], b[16]) ;   // mult.v(2679)
    and (wand_783, a[24], b[15]) ;   // mult.v(2680)
    and (wand_814, a[25], b[14]) ;   // mult.v(2681)
    fa fa_152 (.a(wand_752), .b(wand_783), .cin(wand_814), .s(wfa_s_152), 
       .cout(wfa_cout_152));   // mult.v(2682)
    and (wand_319, a[9], b[31]) ;   // mult.v(2683)
    and (wand_350, a[10], b[30]) ;   // mult.v(2684)
    and (wand_381, a[11], b[29]) ;   // mult.v(2685)
    fa fa_153 (.a(wand_319), .b(wand_350), .cin(wand_381), .s(wfa_s_153), 
       .cout(wfa_cout_153));   // mult.v(2686)
    and (wand_412, a[12], b[28]) ;   // mult.v(2687)
    and (wand_443, a[13], b[27]) ;   // mult.v(2688)
    and (wand_474, a[14], b[26]) ;   // mult.v(2689)
    fa fa_154 (.a(wand_412), .b(wand_443), .cin(wand_474), .s(wfa_s_154), 
       .cout(wfa_cout_154));   // mult.v(2690)
    and (wand_505, a[15], b[25]) ;   // mult.v(2691)
    and (wand_536, a[16], b[24]) ;   // mult.v(2692)
    and (wand_567, a[17], b[23]) ;   // mult.v(2693)
    fa fa_155 (.a(wand_505), .b(wand_536), .cin(wand_567), .s(wfa_s_155), 
       .cout(wfa_cout_155));   // mult.v(2694)
    and (wand_598, a[18], b[22]) ;   // mult.v(2695)
    and (wand_629, a[19], b[21]) ;   // mult.v(2696)
    and (wand_660, a[20], b[20]) ;   // mult.v(2697)
    fa fa_156 (.a(wand_598), .b(wand_629), .cin(wand_660), .s(wfa_s_156), 
       .cout(wfa_cout_156));   // mult.v(2698)
    and (wand_691, a[21], b[19]) ;   // mult.v(2699)
    and (wand_722, a[22], b[18]) ;   // mult.v(2700)
    and (wand_753, a[23], b[17]) ;   // mult.v(2701)
    fa fa_157 (.a(wand_691), .b(wand_722), .cin(wand_753), .s(wfa_s_157), 
       .cout(wfa_cout_157));   // mult.v(2702)
    and (wand_351, a[10], b[31]) ;   // mult.v(2703)
    and (wand_382, a[11], b[30]) ;   // mult.v(2704)
    and (wand_413, a[12], b[29]) ;   // mult.v(2705)
    fa fa_158 (.a(wand_351), .b(wand_382), .cin(wand_413), .s(wfa_s_158), 
       .cout(wfa_cout_158));   // mult.v(2706)
    and (wand_444, a[13], b[28]) ;   // mult.v(2707)
    and (wand_475, a[14], b[27]) ;   // mult.v(2708)
    and (wand_506, a[15], b[26]) ;   // mult.v(2709)
    fa fa_159 (.a(wand_444), .b(wand_475), .cin(wand_506), .s(wfa_s_159), 
       .cout(wfa_cout_159));   // mult.v(2710)
    and (wand_537, a[16], b[25]) ;   // mult.v(2711)
    and (wand_568, a[17], b[24]) ;   // mult.v(2712)
    and (wand_599, a[18], b[23]) ;   // mult.v(2713)
    fa fa_160 (.a(wand_537), .b(wand_568), .cin(wand_599), .s(wfa_s_160), 
       .cout(wfa_cout_160));   // mult.v(2714)
    and (wand_630, a[19], b[22]) ;   // mult.v(2715)
    and (wand_661, a[20], b[21]) ;   // mult.v(2716)
    and (wand_692, a[21], b[20]) ;   // mult.v(2717)
    fa fa_161 (.a(wand_630), .b(wand_661), .cin(wand_692), .s(wfa_s_161), 
       .cout(wfa_cout_161));   // mult.v(2718)
    and (wand_383, a[11], b[31]) ;   // mult.v(2719)
    and (wand_414, a[12], b[30]) ;   // mult.v(2720)
    and (wand_445, a[13], b[29]) ;   // mult.v(2721)
    fa fa_162 (.a(wand_383), .b(wand_414), .cin(wand_445), .s(wfa_s_162), 
       .cout(wfa_cout_162));   // mult.v(2722)
    and (wand_476, a[14], b[28]) ;   // mult.v(2723)
    and (wand_507, a[15], b[27]) ;   // mult.v(2724)
    and (wand_538, a[16], b[26]) ;   // mult.v(2725)
    fa fa_163 (.a(wand_476), .b(wand_507), .cin(wand_538), .s(wfa_s_163), 
       .cout(wfa_cout_163));   // mult.v(2726)
    and (wand_569, a[17], b[25]) ;   // mult.v(2727)
    and (wand_600, a[18], b[24]) ;   // mult.v(2728)
    and (wand_631, a[19], b[23]) ;   // mult.v(2729)
    fa fa_164 (.a(wand_569), .b(wand_600), .cin(wand_631), .s(wfa_s_164), 
       .cout(wfa_cout_164));   // mult.v(2730)
    and (wand_415, a[12], b[31]) ;   // mult.v(2731)
    and (wand_446, a[13], b[30]) ;   // mult.v(2732)
    and (wand_477, a[14], b[29]) ;   // mult.v(2733)
    fa fa_165 (.a(wand_415), .b(wand_446), .cin(wand_477), .s(wfa_s_165), 
       .cout(wfa_cout_165));   // mult.v(2734)
    and (wand_508, a[15], b[28]) ;   // mult.v(2735)
    and (wand_539, a[16], b[27]) ;   // mult.v(2736)
    and (wand_570, a[17], b[26]) ;   // mult.v(2737)
    fa fa_166 (.a(wand_508), .b(wand_539), .cin(wand_570), .s(wfa_s_166), 
       .cout(wfa_cout_166));   // mult.v(2738)
    and (wand_447, a[13], b[31]) ;   // mult.v(2739)
    and (wand_478, a[14], b[30]) ;   // mult.v(2740)
    and (wand_509, a[15], b[29]) ;   // mult.v(2741)
    fa fa_167 (.a(wand_447), .b(wand_478), .cin(wand_509), .s(wfa_s_167), 
       .cout(wfa_cout_167));   // mult.v(2742)
    and (wand_13, a[0], b[13]) ;   // mult.v(2743)
    and (wand_44, a[1], b[12]) ;   // mult.v(2744)
    ha ha_14 (.a(wand_13), .b(wand_44), .s(wha_s_14), .c(wha_c_14));   // mult.v(2745)
    and (wand_14, a[0], b[14]) ;   // mult.v(2746)
    and (wand_45, a[1], b[13]) ;   // mult.v(2747)
    and (wand_76, a[2], b[12]) ;   // mult.v(2748)
    fa fa_168 (.a(wand_14), .b(wand_45), .cin(wand_76), .s(wfa_s_168), 
       .cout(wfa_cout_168));   // mult.v(2749)
    and (wand_107, a[3], b[11]) ;   // mult.v(2750)
    and (wand_138, a[4], b[10]) ;   // mult.v(2751)
    ha ha_15 (.a(wand_107), .b(wand_138), .s(wha_s_15), .c(wha_c_15));   // mult.v(2752)
    and (wand_15, a[0], b[15]) ;   // mult.v(2753)
    and (wand_46, a[1], b[14]) ;   // mult.v(2754)
    and (wand_77, a[2], b[13]) ;   // mult.v(2755)
    fa fa_169 (.a(wand_15), .b(wand_46), .cin(wand_77), .s(wfa_s_169), 
       .cout(wfa_cout_169));   // mult.v(2756)
    and (wand_108, a[3], b[12]) ;   // mult.v(2757)
    and (wand_139, a[4], b[11]) ;   // mult.v(2758)
    and (wand_170, a[5], b[10]) ;   // mult.v(2759)
    fa fa_170 (.a(wand_108), .b(wand_139), .cin(wand_170), .s(wfa_s_170), 
       .cout(wfa_cout_170));   // mult.v(2760)
    and (wand_201, a[6], b[9]) ;   // mult.v(2761)
    and (wand_232, a[7], b[8]) ;   // mult.v(2762)
    ha ha_16 (.a(wand_201), .b(wand_232), .s(wha_s_16), .c(wha_c_16));   // mult.v(2763)
    and (wand_16, a[0], b[16]) ;   // mult.v(2764)
    and (wand_47, a[1], b[15]) ;   // mult.v(2765)
    and (wand_78, a[2], b[14]) ;   // mult.v(2766)
    fa fa_171 (.a(wand_16), .b(wand_47), .cin(wand_78), .s(wfa_s_171), 
       .cout(wfa_cout_171));   // mult.v(2767)
    and (wand_109, a[3], b[13]) ;   // mult.v(2768)
    and (wand_140, a[4], b[12]) ;   // mult.v(2769)
    and (wand_171, a[5], b[11]) ;   // mult.v(2770)
    fa fa_172 (.a(wand_109), .b(wand_140), .cin(wand_171), .s(wfa_s_172), 
       .cout(wfa_cout_172));   // mult.v(2771)
    and (wand_202, a[6], b[10]) ;   // mult.v(2772)
    and (wand_233, a[7], b[9]) ;   // mult.v(2773)
    and (wand_264, a[8], b[8]) ;   // mult.v(2774)
    fa fa_173 (.a(wand_202), .b(wand_233), .cin(wand_264), .s(wfa_s_173), 
       .cout(wfa_cout_173));   // mult.v(2775)
    and (wand_295, a[9], b[7]) ;   // mult.v(2776)
    and (wand_326, a[10], b[6]) ;   // mult.v(2777)
    ha ha_17 (.a(wand_295), .b(wand_326), .s(wha_s_17), .c(wha_c_17));   // mult.v(2778)
    and (wand_17, a[0], b[17]) ;   // mult.v(2779)
    and (wand_48, a[1], b[16]) ;   // mult.v(2780)
    and (wand_79, a[2], b[15]) ;   // mult.v(2781)
    fa fa_174 (.a(wand_17), .b(wand_48), .cin(wand_79), .s(wfa_s_174), 
       .cout(wfa_cout_174));   // mult.v(2782)
    and (wand_110, a[3], b[14]) ;   // mult.v(2783)
    and (wand_141, a[4], b[13]) ;   // mult.v(2784)
    and (wand_172, a[5], b[12]) ;   // mult.v(2785)
    fa fa_175 (.a(wand_110), .b(wand_141), .cin(wand_172), .s(wfa_s_175), 
       .cout(wfa_cout_175));   // mult.v(2786)
    and (wand_203, a[6], b[11]) ;   // mult.v(2787)
    and (wand_234, a[7], b[10]) ;   // mult.v(2788)
    and (wand_265, a[8], b[9]) ;   // mult.v(2789)
    fa fa_176 (.a(wand_203), .b(wand_234), .cin(wand_265), .s(wfa_s_176), 
       .cout(wfa_cout_176));   // mult.v(2790)
    and (wand_296, a[9], b[8]) ;   // mult.v(2791)
    and (wand_327, a[10], b[7]) ;   // mult.v(2792)
    and (wand_358, a[11], b[6]) ;   // mult.v(2793)
    fa fa_177 (.a(wand_296), .b(wand_327), .cin(wand_358), .s(wfa_s_177), 
       .cout(wfa_cout_177));   // mult.v(2794)
    and (wand_389, a[12], b[5]) ;   // mult.v(2795)
    and (wand_420, a[13], b[4]) ;   // mult.v(2796)
    ha ha_18 (.a(wand_389), .b(wand_420), .s(wha_s_18), .c(wha_c_18));   // mult.v(2797)
    and (wand_18, a[0], b[18]) ;   // mult.v(2798)
    and (wand_49, a[1], b[17]) ;   // mult.v(2799)
    and (wand_80, a[2], b[16]) ;   // mult.v(2800)
    fa fa_178 (.a(wand_18), .b(wand_49), .cin(wand_80), .s(wfa_s_178), 
       .cout(wfa_cout_178));   // mult.v(2801)
    and (wand_111, a[3], b[15]) ;   // mult.v(2802)
    and (wand_142, a[4], b[14]) ;   // mult.v(2803)
    and (wand_173, a[5], b[13]) ;   // mult.v(2804)
    fa fa_179 (.a(wand_111), .b(wand_142), .cin(wand_173), .s(wfa_s_179), 
       .cout(wfa_cout_179));   // mult.v(2805)
    and (wand_204, a[6], b[12]) ;   // mult.v(2806)
    and (wand_235, a[7], b[11]) ;   // mult.v(2807)
    and (wand_266, a[8], b[10]) ;   // mult.v(2808)
    fa fa_180 (.a(wand_204), .b(wand_235), .cin(wand_266), .s(wfa_s_180), 
       .cout(wfa_cout_180));   // mult.v(2809)
    and (wand_297, a[9], b[9]) ;   // mult.v(2810)
    and (wand_328, a[10], b[8]) ;   // mult.v(2811)
    and (wand_359, a[11], b[7]) ;   // mult.v(2812)
    fa fa_181 (.a(wand_297), .b(wand_328), .cin(wand_359), .s(wfa_s_181), 
       .cout(wfa_cout_181));   // mult.v(2813)
    and (wand_390, a[12], b[6]) ;   // mult.v(2814)
    and (wand_421, a[13], b[5]) ;   // mult.v(2815)
    and (wand_452, a[14], b[4]) ;   // mult.v(2816)
    fa fa_182 (.a(wand_390), .b(wand_421), .cin(wand_452), .s(wfa_s_182), 
       .cout(wfa_cout_182));   // mult.v(2817)
    and (wand_483, a[15], b[3]) ;   // mult.v(2818)
    and (wand_514, a[16], b[2]) ;   // mult.v(2819)
    ha ha_19 (.a(wand_483), .b(wand_514), .s(wha_s_19), .c(wha_c_19));   // mult.v(2820)
    and (wand_81, a[2], b[17]) ;   // mult.v(2821)
    and (wand_112, a[3], b[16]) ;   // mult.v(2822)
    and (wand_143, a[4], b[15]) ;   // mult.v(2823)
    fa fa_183 (.a(wand_81), .b(wand_112), .cin(wand_143), .s(wfa_s_183), 
       .cout(wfa_cout_183));   // mult.v(2824)
    and (wand_174, a[5], b[14]) ;   // mult.v(2825)
    and (wand_205, a[6], b[13]) ;   // mult.v(2826)
    and (wand_236, a[7], b[12]) ;   // mult.v(2827)
    fa fa_184 (.a(wand_174), .b(wand_205), .cin(wand_236), .s(wfa_s_184), 
       .cout(wfa_cout_184));   // mult.v(2828)
    and (wand_267, a[8], b[11]) ;   // mult.v(2829)
    and (wand_298, a[9], b[10]) ;   // mult.v(2830)
    and (wand_329, a[10], b[9]) ;   // mult.v(2831)
    fa fa_185 (.a(wand_267), .b(wand_298), .cin(wand_329), .s(wfa_s_185), 
       .cout(wfa_cout_185));   // mult.v(2832)
    and (wand_360, a[11], b[8]) ;   // mult.v(2833)
    and (wand_391, a[12], b[7]) ;   // mult.v(2834)
    and (wand_422, a[13], b[6]) ;   // mult.v(2835)
    fa fa_186 (.a(wand_360), .b(wand_391), .cin(wand_422), .s(wfa_s_186), 
       .cout(wfa_cout_186));   // mult.v(2836)
    and (wand_453, a[14], b[5]) ;   // mult.v(2837)
    and (wand_484, a[15], b[4]) ;   // mult.v(2838)
    and (wand_515, a[16], b[3]) ;   // mult.v(2839)
    fa fa_187 (.a(wand_453), .b(wand_484), .cin(wand_515), .s(wfa_s_187), 
       .cout(wfa_cout_187));   // mult.v(2840)
    and (wand_546, a[17], b[2]) ;   // mult.v(2841)
    and (wand_577, a[18], b[1]) ;   // mult.v(2842)
    and (wand_608, a[19], b[0]) ;   // mult.v(2843)
    fa fa_188 (.a(wand_546), .b(wand_577), .cin(wand_608), .s(wfa_s_188), 
       .cout(wfa_cout_188));   // mult.v(2844)
    and (wand_175, a[5], b[15]) ;   // mult.v(2845)
    and (wand_206, a[6], b[14]) ;   // mult.v(2846)
    and (wand_237, a[7], b[13]) ;   // mult.v(2847)
    fa fa_189 (.a(wand_175), .b(wand_206), .cin(wand_237), .s(wfa_s_189), 
       .cout(wfa_cout_189));   // mult.v(2848)
    and (wand_268, a[8], b[12]) ;   // mult.v(2849)
    and (wand_299, a[9], b[11]) ;   // mult.v(2850)
    and (wand_330, a[10], b[10]) ;   // mult.v(2851)
    fa fa_190 (.a(wand_268), .b(wand_299), .cin(wand_330), .s(wfa_s_190), 
       .cout(wfa_cout_190));   // mult.v(2852)
    and (wand_361, a[11], b[9]) ;   // mult.v(2853)
    and (wand_392, a[12], b[8]) ;   // mult.v(2854)
    and (wand_423, a[13], b[7]) ;   // mult.v(2855)
    fa fa_191 (.a(wand_361), .b(wand_392), .cin(wand_423), .s(wfa_s_191), 
       .cout(wfa_cout_191));   // mult.v(2856)
    and (wand_454, a[14], b[6]) ;   // mult.v(2857)
    and (wand_485, a[15], b[5]) ;   // mult.v(2858)
    and (wand_516, a[16], b[4]) ;   // mult.v(2859)
    fa fa_192 (.a(wand_454), .b(wand_485), .cin(wand_516), .s(wfa_s_192), 
       .cout(wfa_cout_192));   // mult.v(2860)
    and (wand_547, a[17], b[3]) ;   // mult.v(2861)
    and (wand_578, a[18], b[2]) ;   // mult.v(2862)
    and (wand_609, a[19], b[1]) ;   // mult.v(2863)
    fa fa_193 (.a(wand_547), .b(wand_578), .cin(wand_609), .s(wfa_s_193), 
       .cout(wfa_cout_193));   // mult.v(2864)
    and (wand_640, a[20], b[0]) ;   // mult.v(2865)
    fa fa_194 (.a(wand_640), .b(wha_c_5), .cin(wfa_s_15), .s(wfa_s_194), 
       .cout(wfa_cout_194));   // mult.v(2866)
    and (wand_269, a[8], b[13]) ;   // mult.v(2867)
    and (wand_300, a[9], b[12]) ;   // mult.v(2868)
    and (wand_331, a[10], b[11]) ;   // mult.v(2869)
    fa fa_195 (.a(wand_269), .b(wand_300), .cin(wand_331), .s(wfa_s_195), 
       .cout(wfa_cout_195));   // mult.v(2870)
    and (wand_362, a[11], b[10]) ;   // mult.v(2871)
    and (wand_393, a[12], b[9]) ;   // mult.v(2872)
    and (wand_424, a[13], b[8]) ;   // mult.v(2873)
    fa fa_196 (.a(wand_362), .b(wand_393), .cin(wand_424), .s(wfa_s_196), 
       .cout(wfa_cout_196));   // mult.v(2874)
    and (wand_455, a[14], b[7]) ;   // mult.v(2875)
    and (wand_486, a[15], b[6]) ;   // mult.v(2876)
    and (wand_517, a[16], b[5]) ;   // mult.v(2877)
    fa fa_197 (.a(wand_455), .b(wand_486), .cin(wand_517), .s(wfa_s_197), 
       .cout(wfa_cout_197));   // mult.v(2878)
    and (wand_548, a[17], b[4]) ;   // mult.v(2879)
    and (wand_579, a[18], b[3]) ;   // mult.v(2880)
    and (wand_610, a[19], b[2]) ;   // mult.v(2881)
    fa fa_198 (.a(wand_548), .b(wand_579), .cin(wand_610), .s(wfa_s_198), 
       .cout(wfa_cout_198));   // mult.v(2882)
    and (wand_641, a[20], b[1]) ;   // mult.v(2883)
    and (wand_672, a[21], b[0]) ;   // mult.v(2884)
    fa fa_199 (.a(wand_641), .b(wand_672), .cin(wfa_cout_15), .s(wfa_s_199), 
       .cout(wfa_cout_199));   // mult.v(2885)
    fa fa_200 (.a(wha_c_6), .b(wfa_s_16), .cin(wfa_s_17), .s(wfa_s_200), 
       .cout(wfa_cout_200));   // mult.v(2886)
    and (wand_363, a[11], b[11]) ;   // mult.v(2887)
    and (wand_394, a[12], b[10]) ;   // mult.v(2888)
    and (wand_425, a[13], b[9]) ;   // mult.v(2889)
    fa fa_201 (.a(wand_363), .b(wand_394), .cin(wand_425), .s(wfa_s_201), 
       .cout(wfa_cout_201));   // mult.v(2890)
    and (wand_456, a[14], b[8]) ;   // mult.v(2891)
    and (wand_487, a[15], b[7]) ;   // mult.v(2892)
    and (wand_518, a[16], b[6]) ;   // mult.v(2893)
    fa fa_202 (.a(wand_456), .b(wand_487), .cin(wand_518), .s(wfa_s_202), 
       .cout(wfa_cout_202));   // mult.v(2894)
    and (wand_549, a[17], b[5]) ;   // mult.v(2895)
    and (wand_580, a[18], b[4]) ;   // mult.v(2896)
    and (wand_611, a[19], b[3]) ;   // mult.v(2897)
    fa fa_203 (.a(wand_549), .b(wand_580), .cin(wand_611), .s(wfa_s_203), 
       .cout(wfa_cout_203));   // mult.v(2898)
    and (wand_642, a[20], b[2]) ;   // mult.v(2899)
    and (wand_673, a[21], b[1]) ;   // mult.v(2900)
    and (wand_704, a[22], b[0]) ;   // mult.v(2901)
    fa fa_204 (.a(wand_642), .b(wand_673), .cin(wand_704), .s(wfa_s_204), 
       .cout(wfa_cout_204));   // mult.v(2902)
    fa fa_205 (.a(wfa_cout_16), .b(wfa_cout_17), .cin(wha_c_7), .s(wfa_s_205), 
       .cout(wfa_cout_205));   // mult.v(2903)
    fa fa_206 (.a(wfa_s_18), .b(wfa_s_19), .cin(wfa_s_20), .s(wfa_s_206), 
       .cout(wfa_cout_206));   // mult.v(2904)
    and (wand_457, a[14], b[9]) ;   // mult.v(2905)
    and (wand_488, a[15], b[8]) ;   // mult.v(2906)
    and (wand_519, a[16], b[7]) ;   // mult.v(2907)
    fa fa_207 (.a(wand_457), .b(wand_488), .cin(wand_519), .s(wfa_s_207), 
       .cout(wfa_cout_207));   // mult.v(2908)
    and (wand_550, a[17], b[6]) ;   // mult.v(2909)
    and (wand_581, a[18], b[5]) ;   // mult.v(2910)
    and (wand_612, a[19], b[4]) ;   // mult.v(2911)
    fa fa_208 (.a(wand_550), .b(wand_581), .cin(wand_612), .s(wfa_s_208), 
       .cout(wfa_cout_208));   // mult.v(2912)
    and (wand_643, a[20], b[3]) ;   // mult.v(2913)
    and (wand_674, a[21], b[2]) ;   // mult.v(2914)
    and (wand_705, a[22], b[1]) ;   // mult.v(2915)
    fa fa_209 (.a(wand_643), .b(wand_674), .cin(wand_705), .s(wfa_s_209), 
       .cout(wfa_cout_209));   // mult.v(2916)
    and (wand_736, a[23], b[0]) ;   // mult.v(2917)
    fa fa_210 (.a(wand_736), .b(wfa_cout_18), .cin(wfa_cout_19), .s(wfa_s_210), 
       .cout(wfa_cout_210));   // mult.v(2918)
    fa fa_211 (.a(wfa_cout_20), .b(wha_c_8), .cin(wfa_s_21), .s(wfa_s_211), 
       .cout(wfa_cout_211));   // mult.v(2919)
    fa fa_212 (.a(wfa_s_22), .b(wfa_s_23), .cin(wfa_s_24), .s(wfa_s_212), 
       .cout(wfa_cout_212));   // mult.v(2920)
    and (wand_551, a[17], b[7]) ;   // mult.v(2921)
    and (wand_582, a[18], b[6]) ;   // mult.v(2922)
    and (wand_613, a[19], b[5]) ;   // mult.v(2923)
    fa fa_213 (.a(wand_551), .b(wand_582), .cin(wand_613), .s(wfa_s_213), 
       .cout(wfa_cout_213));   // mult.v(2924)
    and (wand_644, a[20], b[4]) ;   // mult.v(2925)
    and (wand_675, a[21], b[3]) ;   // mult.v(2926)
    and (wand_706, a[22], b[2]) ;   // mult.v(2927)
    fa fa_214 (.a(wand_644), .b(wand_675), .cin(wand_706), .s(wfa_s_214), 
       .cout(wfa_cout_214));   // mult.v(2928)
    and (wand_737, a[23], b[1]) ;   // mult.v(2929)
    and (wand_768, a[24], b[0]) ;   // mult.v(2930)
    fa fa_215 (.a(wand_737), .b(wand_768), .cin(wfa_cout_21), .s(wfa_s_215), 
       .cout(wfa_cout_215));   // mult.v(2931)
    fa fa_216 (.a(wfa_cout_22), .b(wfa_cout_23), .cin(wfa_cout_24), .s(wfa_s_216), 
       .cout(wfa_cout_216));   // mult.v(2932)
    fa fa_217 (.a(wha_c_9), .b(wfa_s_25), .cin(wfa_s_26), .s(wfa_s_217), 
       .cout(wfa_cout_217));   // mult.v(2933)
    fa fa_218 (.a(wfa_s_27), .b(wfa_s_28), .cin(wfa_s_29), .s(wfa_s_218), 
       .cout(wfa_cout_218));   // mult.v(2934)
    and (wand_645, a[20], b[5]) ;   // mult.v(2935)
    and (wand_676, a[21], b[4]) ;   // mult.v(2936)
    and (wand_707, a[22], b[3]) ;   // mult.v(2937)
    fa fa_219 (.a(wand_645), .b(wand_676), .cin(wand_707), .s(wfa_s_219), 
       .cout(wfa_cout_219));   // mult.v(2938)
    and (wand_738, a[23], b[2]) ;   // mult.v(2939)
    and (wand_769, a[24], b[1]) ;   // mult.v(2940)
    and (wand_800, a[25], b[0]) ;   // mult.v(2941)
    fa fa_220 (.a(wand_738), .b(wand_769), .cin(wand_800), .s(wfa_s_220), 
       .cout(wfa_cout_220));   // mult.v(2942)
    fa fa_221 (.a(wfa_cout_25), .b(wfa_cout_26), .cin(wfa_cout_27), .s(wfa_s_221), 
       .cout(wfa_cout_221));   // mult.v(2943)
    fa fa_222 (.a(wfa_cout_28), .b(wfa_cout_29), .cin(wha_c_10), .s(wfa_s_222), 
       .cout(wfa_cout_222));   // mult.v(2944)
    fa fa_223 (.a(wfa_s_30), .b(wfa_s_31), .cin(wfa_s_32), .s(wfa_s_223), 
       .cout(wfa_cout_223));   // mult.v(2945)
    fa fa_224 (.a(wfa_s_33), .b(wfa_s_34), .cin(wfa_s_35), .s(wfa_s_224), 
       .cout(wfa_cout_224));   // mult.v(2946)
    and (wand_739, a[23], b[3]) ;   // mult.v(2947)
    and (wand_770, a[24], b[2]) ;   // mult.v(2948)
    and (wand_801, a[25], b[1]) ;   // mult.v(2949)
    fa fa_225 (.a(wand_739), .b(wand_770), .cin(wand_801), .s(wfa_s_225), 
       .cout(wfa_cout_225));   // mult.v(2950)
    and (wand_832, a[26], b[0]) ;   // mult.v(2951)
    fa fa_226 (.a(wand_832), .b(wfa_cout_30), .cin(wfa_cout_31), .s(wfa_s_226), 
       .cout(wfa_cout_226));   // mult.v(2952)
    fa fa_227 (.a(wfa_cout_32), .b(wfa_cout_33), .cin(wfa_cout_34), .s(wfa_s_227), 
       .cout(wfa_cout_227));   // mult.v(2953)
    fa fa_228 (.a(wfa_cout_35), .b(wha_c_11), .cin(wfa_s_36), .s(wfa_s_228), 
       .cout(wfa_cout_228));   // mult.v(2954)
    fa fa_229 (.a(wfa_s_37), .b(wfa_s_38), .cin(wfa_s_39), .s(wfa_s_229), 
       .cout(wfa_cout_229));   // mult.v(2955)
    fa fa_230 (.a(wfa_s_40), .b(wfa_s_41), .cin(wfa_s_42), .s(wfa_s_230), 
       .cout(wfa_cout_230));   // mult.v(2956)
    and (wand_833, a[26], b[1]) ;   // mult.v(2957)
    and (wand_864, a[27], b[0]) ;   // mult.v(2958)
    fa fa_231 (.a(wand_833), .b(wand_864), .cin(wfa_cout_36), .s(wfa_s_231), 
       .cout(wfa_cout_231));   // mult.v(2959)
    fa fa_232 (.a(wfa_cout_37), .b(wfa_cout_38), .cin(wfa_cout_39), .s(wfa_s_232), 
       .cout(wfa_cout_232));   // mult.v(2960)
    fa fa_233 (.a(wfa_cout_40), .b(wfa_cout_41), .cin(wfa_cout_42), .s(wfa_s_233), 
       .cout(wfa_cout_233));   // mult.v(2961)
    fa fa_234 (.a(wha_c_12), .b(wfa_s_43), .cin(wfa_s_44), .s(wfa_s_234), 
       .cout(wfa_cout_234));   // mult.v(2962)
    fa fa_235 (.a(wfa_s_45), .b(wfa_s_46), .cin(wfa_s_47), .s(wfa_s_235), 
       .cout(wfa_cout_235));   // mult.v(2963)
    fa fa_236 (.a(wfa_s_48), .b(wfa_s_49), .cin(wfa_s_50), .s(wfa_s_236), 
       .cout(wfa_cout_236));   // mult.v(2964)
    fa fa_237 (.a(wha_s_0), .b(wfa_cout_43), .cin(wfa_cout_44), .s(wfa_s_237), 
       .cout(wfa_cout_237));   // mult.v(2965)
    fa fa_238 (.a(wfa_cout_45), .b(wfa_cout_46), .cin(wfa_cout_47), .s(wfa_s_238), 
       .cout(wfa_cout_238));   // mult.v(2966)
    fa fa_239 (.a(wfa_cout_48), .b(wfa_cout_49), .cin(wfa_cout_50), .s(wfa_s_239), 
       .cout(wfa_cout_239));   // mult.v(2967)
    fa fa_240 (.a(wha_c_13), .b(wfa_s_51), .cin(wfa_s_52), .s(wfa_s_240), 
       .cout(wfa_cout_240));   // mult.v(2968)
    fa fa_241 (.a(wfa_s_53), .b(wfa_s_54), .cin(wfa_s_55), .s(wfa_s_241), 
       .cout(wfa_cout_241));   // mult.v(2969)
    fa fa_242 (.a(wfa_s_56), .b(wfa_s_57), .cin(wfa_s_58), .s(wfa_s_242), 
       .cout(wfa_cout_242));   // mult.v(2970)
    fa fa_243 (.a(wha_s_1), .b(wfa_cout_51), .cin(wfa_cout_52), .s(wfa_s_243), 
       .cout(wfa_cout_243));   // mult.v(2971)
    fa fa_244 (.a(wfa_cout_53), .b(wfa_cout_54), .cin(wfa_cout_55), .s(wfa_s_244), 
       .cout(wfa_cout_244));   // mult.v(2972)
    fa fa_245 (.a(wfa_cout_56), .b(wfa_cout_57), .cin(wfa_cout_58), .s(wfa_s_245), 
       .cout(wfa_cout_245));   // mult.v(2973)
    fa fa_246 (.a(wfa_cout_59), .b(wfa_s_60), .cin(wfa_s_61), .s(wfa_s_246), 
       .cout(wfa_cout_246));   // mult.v(2974)
    fa fa_247 (.a(wfa_s_62), .b(wfa_s_63), .cin(wfa_s_64), .s(wfa_s_247), 
       .cout(wfa_cout_247));   // mult.v(2975)
    fa fa_248 (.a(wfa_s_65), .b(wfa_s_66), .cin(wfa_s_67), .s(wfa_s_248), 
       .cout(wfa_cout_248));   // mult.v(2976)
    fa fa_249 (.a(wha_s_2), .b(wfa_cout_60), .cin(wfa_cout_61), .s(wfa_s_249), 
       .cout(wfa_cout_249));   // mult.v(2977)
    fa fa_250 (.a(wfa_cout_62), .b(wfa_cout_63), .cin(wfa_cout_64), .s(wfa_s_250), 
       .cout(wfa_cout_250));   // mult.v(2978)
    fa fa_251 (.a(wfa_cout_65), .b(wfa_cout_66), .cin(wfa_cout_67), .s(wfa_s_251), 
       .cout(wfa_cout_251));   // mult.v(2979)
    fa fa_252 (.a(wfa_cout_68), .b(wfa_s_69), .cin(wfa_s_70), .s(wfa_s_252), 
       .cout(wfa_cout_252));   // mult.v(2980)
    fa fa_253 (.a(wfa_s_71), .b(wfa_s_72), .cin(wfa_s_73), .s(wfa_s_253), 
       .cout(wfa_cout_253));   // mult.v(2981)
    fa fa_254 (.a(wfa_s_74), .b(wfa_s_75), .cin(wfa_s_76), .s(wfa_s_254), 
       .cout(wfa_cout_254));   // mult.v(2982)
    fa fa_255 (.a(wha_s_3), .b(wfa_cout_69), .cin(wfa_cout_70), .s(wfa_s_255), 
       .cout(wfa_cout_255));   // mult.v(2983)
    fa fa_256 (.a(wfa_cout_71), .b(wfa_cout_72), .cin(wfa_cout_73), .s(wfa_s_256), 
       .cout(wfa_cout_256));   // mult.v(2984)
    fa fa_257 (.a(wfa_cout_74), .b(wfa_cout_75), .cin(wfa_cout_76), .s(wfa_s_257), 
       .cout(wfa_cout_257));   // mult.v(2985)
    fa fa_258 (.a(wfa_cout_77), .b(wfa_s_78), .cin(wfa_s_79), .s(wfa_s_258), 
       .cout(wfa_cout_258));   // mult.v(2986)
    fa fa_259 (.a(wfa_s_80), .b(wfa_s_81), .cin(wfa_s_82), .s(wfa_s_259), 
       .cout(wfa_cout_259));   // mult.v(2987)
    fa fa_260 (.a(wfa_s_83), .b(wfa_s_84), .cin(wfa_s_85), .s(wfa_s_260), 
       .cout(wfa_cout_260));   // mult.v(2988)
    fa fa_261 (.a(wha_s_4), .b(wfa_cout_78), .cin(wfa_cout_79), .s(wfa_s_261), 
       .cout(wfa_cout_261));   // mult.v(2989)
    fa fa_262 (.a(wfa_cout_80), .b(wfa_cout_81), .cin(wfa_cout_82), .s(wfa_s_262), 
       .cout(wfa_cout_262));   // mult.v(2990)
    fa fa_263 (.a(wfa_cout_83), .b(wfa_cout_84), .cin(wfa_cout_85), .s(wfa_s_263), 
       .cout(wfa_cout_263));   // mult.v(2991)
    fa fa_264 (.a(wfa_cout_86), .b(wfa_s_87), .cin(wfa_s_88), .s(wfa_s_264), 
       .cout(wfa_cout_264));   // mult.v(2992)
    fa fa_265 (.a(wfa_s_89), .b(wfa_s_90), .cin(wfa_s_91), .s(wfa_s_265), 
       .cout(wfa_cout_265));   // mult.v(2993)
    fa fa_266 (.a(wfa_s_92), .b(wfa_s_93), .cin(wfa_s_94), .s(wfa_s_266), 
       .cout(wfa_cout_266));   // mult.v(2994)
    fa fa_267 (.a(wfa_s_11), .b(wfa_cout_87), .cin(wfa_cout_88), .s(wfa_s_267), 
       .cout(wfa_cout_267));   // mult.v(2995)
    fa fa_268 (.a(wfa_cout_89), .b(wfa_cout_90), .cin(wfa_cout_91), .s(wfa_s_268), 
       .cout(wfa_cout_268));   // mult.v(2996)
    fa fa_269 (.a(wfa_cout_92), .b(wfa_cout_93), .cin(wfa_cout_94), .s(wfa_s_269), 
       .cout(wfa_cout_269));   // mult.v(2997)
    fa fa_270 (.a(wfa_cout_95), .b(wfa_s_96), .cin(wfa_s_97), .s(wfa_s_270), 
       .cout(wfa_cout_270));   // mult.v(2998)
    fa fa_271 (.a(wfa_s_98), .b(wfa_s_99), .cin(wfa_s_100), .s(wfa_s_271), 
       .cout(wfa_cout_271));   // mult.v(2999)
    fa fa_272 (.a(wfa_s_101), .b(wfa_s_102), .cin(wfa_s_103), .s(wfa_s_272), 
       .cout(wfa_cout_272));   // mult.v(3000)
    fa fa_273 (.a(wfa_s_13), .b(wfa_cout_96), .cin(wfa_cout_97), .s(wfa_s_273), 
       .cout(wfa_cout_273));   // mult.v(3001)
    fa fa_274 (.a(wfa_cout_98), .b(wfa_cout_99), .cin(wfa_cout_100), .s(wfa_s_274), 
       .cout(wfa_cout_274));   // mult.v(3002)
    fa fa_275 (.a(wfa_cout_101), .b(wfa_cout_102), .cin(wfa_cout_103), 
       .s(wfa_s_275), .cout(wfa_cout_275));   // mult.v(3003)
    fa fa_276 (.a(wfa_cout_104), .b(wfa_s_105), .cin(wfa_s_106), .s(wfa_s_276), 
       .cout(wfa_cout_276));   // mult.v(3004)
    fa fa_277 (.a(wfa_s_107), .b(wfa_s_108), .cin(wfa_s_109), .s(wfa_s_277), 
       .cout(wfa_cout_277));   // mult.v(3005)
    fa fa_278 (.a(wfa_s_110), .b(wfa_s_111), .cin(wfa_s_112), .s(wfa_s_278), 
       .cout(wfa_cout_278));   // mult.v(3006)
    fa fa_279 (.a(wfa_s_14), .b(wfa_cout_105), .cin(wfa_cout_106), .s(wfa_s_279), 
       .cout(wfa_cout_279));   // mult.v(3007)
    fa fa_280 (.a(wfa_cout_107), .b(wfa_cout_108), .cin(wfa_cout_109), 
       .s(wfa_s_280), .cout(wfa_cout_280));   // mult.v(3008)
    fa fa_281 (.a(wfa_cout_110), .b(wfa_cout_111), .cin(wfa_cout_112), 
       .s(wfa_s_281), .cout(wfa_cout_281));   // mult.v(3009)
    fa fa_282 (.a(wfa_cout_113), .b(wfa_s_114), .cin(wfa_s_115), .s(wfa_s_282), 
       .cout(wfa_cout_282));   // mult.v(3010)
    fa fa_283 (.a(wfa_s_116), .b(wfa_s_117), .cin(wfa_s_118), .s(wfa_s_283), 
       .cout(wfa_cout_283));   // mult.v(3011)
    fa fa_284 (.a(wfa_s_119), .b(wfa_s_120), .cin(wfa_s_121), .s(wfa_s_284), 
       .cout(wfa_cout_284));   // mult.v(3012)
    fa fa_285 (.a(wfa_cout_14), .b(wfa_cout_114), .cin(wfa_cout_115), 
       .s(wfa_s_285), .cout(wfa_cout_285));   // mult.v(3013)
    fa fa_286 (.a(wfa_cout_116), .b(wfa_cout_117), .cin(wfa_cout_118), 
       .s(wfa_s_286), .cout(wfa_cout_286));   // mult.v(3014)
    fa fa_287 (.a(wfa_cout_119), .b(wfa_cout_120), .cin(wfa_cout_121), 
       .s(wfa_s_287), .cout(wfa_cout_287));   // mult.v(3015)
    fa fa_288 (.a(wfa_cout_122), .b(wfa_s_123), .cin(wfa_s_124), .s(wfa_s_288), 
       .cout(wfa_cout_288));   // mult.v(3016)
    fa fa_289 (.a(wfa_s_125), .b(wfa_s_126), .cin(wfa_s_127), .s(wfa_s_289), 
       .cout(wfa_cout_289));   // mult.v(3017)
    fa fa_290 (.a(wfa_s_128), .b(wfa_s_129), .cin(wfa_s_130), .s(wfa_s_290), 
       .cout(wfa_cout_290));   // mult.v(3018)
    and (wand_967, a[30], b[7]) ;   // mult.v(3019)
    and (wand_998, a[31], b[6]) ;   // mult.v(3020)
    fa fa_291 (.a(wand_967), .b(wand_998), .cin(wfa_cout_123), .s(wfa_s_291), 
       .cout(wfa_cout_291));   // mult.v(3021)
    fa fa_292 (.a(wfa_cout_124), .b(wfa_cout_125), .cin(wfa_cout_126), 
       .s(wfa_s_292), .cout(wfa_cout_292));   // mult.v(3022)
    fa fa_293 (.a(wfa_cout_127), .b(wfa_cout_128), .cin(wfa_cout_129), 
       .s(wfa_s_293), .cout(wfa_cout_293));   // mult.v(3023)
    fa fa_294 (.a(wfa_cout_130), .b(wfa_cout_131), .cin(wfa_s_132), .s(wfa_s_294), 
       .cout(wfa_cout_294));   // mult.v(3024)
    fa fa_295 (.a(wfa_s_133), .b(wfa_s_134), .cin(wfa_s_135), .s(wfa_s_295), 
       .cout(wfa_cout_295));   // mult.v(3025)
    fa fa_296 (.a(wfa_s_136), .b(wfa_s_137), .cin(wfa_s_138), .s(wfa_s_296), 
       .cout(wfa_cout_296));   // mult.v(3026)
    and (wand_906, a[28], b[10]) ;   // mult.v(3027)
    and (wand_937, a[29], b[9]) ;   // mult.v(3028)
    and (wand_968, a[30], b[8]) ;   // mult.v(3029)
    fa fa_297 (.a(wand_906), .b(wand_937), .cin(wand_968), .s(wfa_s_297), 
       .cout(wfa_cout_297));   // mult.v(3030)
    and (wand_999, a[31], b[7]) ;   // mult.v(3031)
    fa fa_298 (.a(wand_999), .b(wfa_cout_132), .cin(wfa_cout_133), .s(wfa_s_298), 
       .cout(wfa_cout_298));   // mult.v(3032)
    fa fa_299 (.a(wfa_cout_134), .b(wfa_cout_135), .cin(wfa_cout_136), 
       .s(wfa_s_299), .cout(wfa_cout_299));   // mult.v(3033)
    fa fa_300 (.a(wfa_cout_137), .b(wfa_cout_138), .cin(wfa_cout_139), 
       .s(wfa_s_300), .cout(wfa_cout_300));   // mult.v(3034)
    fa fa_301 (.a(wfa_s_140), .b(wfa_s_141), .cin(wfa_s_142), .s(wfa_s_301), 
       .cout(wfa_cout_301));   // mult.v(3035)
    fa fa_302 (.a(wfa_s_143), .b(wfa_s_144), .cin(wfa_s_145), .s(wfa_s_302), 
       .cout(wfa_cout_302));   // mult.v(3036)
    and (wand_845, a[26], b[13]) ;   // mult.v(3037)
    and (wand_876, a[27], b[12]) ;   // mult.v(3038)
    and (wand_907, a[28], b[11]) ;   // mult.v(3039)
    fa fa_303 (.a(wand_845), .b(wand_876), .cin(wand_907), .s(wfa_s_303), 
       .cout(wfa_cout_303));   // mult.v(3040)
    and (wand_938, a[29], b[10]) ;   // mult.v(3041)
    and (wand_969, a[30], b[9]) ;   // mult.v(3042)
    and (wand_1000, a[31], b[8]) ;   // mult.v(3043)
    fa fa_304 (.a(wand_938), .b(wand_969), .cin(wand_1000), .s(wfa_s_304), 
       .cout(wfa_cout_304));   // mult.v(3044)
    fa fa_305 (.a(wfa_cout_140), .b(wfa_cout_141), .cin(wfa_cout_142), 
       .s(wfa_s_305), .cout(wfa_cout_305));   // mult.v(3045)
    fa fa_306 (.a(wfa_cout_143), .b(wfa_cout_144), .cin(wfa_cout_145), 
       .s(wfa_s_306), .cout(wfa_cout_306));   // mult.v(3046)
    fa fa_307 (.a(wfa_cout_146), .b(wfa_s_147), .cin(wfa_s_148), .s(wfa_s_307), 
       .cout(wfa_cout_307));   // mult.v(3047)
    fa fa_308 (.a(wfa_s_149), .b(wfa_s_150), .cin(wfa_s_151), .s(wfa_s_308), 
       .cout(wfa_cout_308));   // mult.v(3048)
    and (wand_784, a[24], b[16]) ;   // mult.v(3049)
    and (wand_815, a[25], b[15]) ;   // mult.v(3050)
    and (wand_846, a[26], b[14]) ;   // mult.v(3051)
    fa fa_309 (.a(wand_784), .b(wand_815), .cin(wand_846), .s(wfa_s_309), 
       .cout(wfa_cout_309));   // mult.v(3052)
    and (wand_877, a[27], b[13]) ;   // mult.v(3053)
    and (wand_908, a[28], b[12]) ;   // mult.v(3054)
    and (wand_939, a[29], b[11]) ;   // mult.v(3055)
    fa fa_310 (.a(wand_877), .b(wand_908), .cin(wand_939), .s(wfa_s_310), 
       .cout(wfa_cout_310));   // mult.v(3056)
    and (wand_970, a[30], b[10]) ;   // mult.v(3057)
    and (wand_1001, a[31], b[9]) ;   // mult.v(3058)
    fa fa_311 (.a(wand_970), .b(wand_1001), .cin(wfa_cout_147), .s(wfa_s_311), 
       .cout(wfa_cout_311));   // mult.v(3059)
    fa fa_312 (.a(wfa_cout_148), .b(wfa_cout_149), .cin(wfa_cout_150), 
       .s(wfa_s_312), .cout(wfa_cout_312));   // mult.v(3060)
    fa fa_313 (.a(wfa_cout_151), .b(wfa_cout_152), .cin(wfa_s_153), .s(wfa_s_313), 
       .cout(wfa_cout_313));   // mult.v(3061)
    fa fa_314 (.a(wfa_s_154), .b(wfa_s_155), .cin(wfa_s_156), .s(wfa_s_314), 
       .cout(wfa_cout_314));   // mult.v(3062)
    and (wand_723, a[22], b[19]) ;   // mult.v(3063)
    and (wand_754, a[23], b[18]) ;   // mult.v(3064)
    and (wand_785, a[24], b[17]) ;   // mult.v(3065)
    fa fa_315 (.a(wand_723), .b(wand_754), .cin(wand_785), .s(wfa_s_315), 
       .cout(wfa_cout_315));   // mult.v(3066)
    and (wand_816, a[25], b[16]) ;   // mult.v(3067)
    and (wand_847, a[26], b[15]) ;   // mult.v(3068)
    and (wand_878, a[27], b[14]) ;   // mult.v(3069)
    fa fa_316 (.a(wand_816), .b(wand_847), .cin(wand_878), .s(wfa_s_316), 
       .cout(wfa_cout_316));   // mult.v(3070)
    and (wand_909, a[28], b[13]) ;   // mult.v(3071)
    and (wand_940, a[29], b[12]) ;   // mult.v(3072)
    and (wand_971, a[30], b[11]) ;   // mult.v(3073)
    fa fa_317 (.a(wand_909), .b(wand_940), .cin(wand_971), .s(wfa_s_317), 
       .cout(wfa_cout_317));   // mult.v(3074)
    and (wand_1002, a[31], b[10]) ;   // mult.v(3075)
    fa fa_318 (.a(wand_1002), .b(wfa_cout_153), .cin(wfa_cout_154), .s(wfa_s_318), 
       .cout(wfa_cout_318));   // mult.v(3076)
    fa fa_319 (.a(wfa_cout_155), .b(wfa_cout_156), .cin(wfa_cout_157), 
       .s(wfa_s_319), .cout(wfa_cout_319));   // mult.v(3077)
    fa fa_320 (.a(wfa_s_158), .b(wfa_s_159), .cin(wfa_s_160), .s(wfa_s_320), 
       .cout(wfa_cout_320));   // mult.v(3078)
    and (wand_662, a[20], b[22]) ;   // mult.v(3079)
    and (wand_693, a[21], b[21]) ;   // mult.v(3080)
    and (wand_724, a[22], b[20]) ;   // mult.v(3081)
    fa fa_321 (.a(wand_662), .b(wand_693), .cin(wand_724), .s(wfa_s_321), 
       .cout(wfa_cout_321));   // mult.v(3082)
    and (wand_755, a[23], b[19]) ;   // mult.v(3083)
    and (wand_786, a[24], b[18]) ;   // mult.v(3084)
    and (wand_817, a[25], b[17]) ;   // mult.v(3085)
    fa fa_322 (.a(wand_755), .b(wand_786), .cin(wand_817), .s(wfa_s_322), 
       .cout(wfa_cout_322));   // mult.v(3086)
    and (wand_848, a[26], b[16]) ;   // mult.v(3087)
    and (wand_879, a[27], b[15]) ;   // mult.v(3088)
    and (wand_910, a[28], b[14]) ;   // mult.v(3089)
    fa fa_323 (.a(wand_848), .b(wand_879), .cin(wand_910), .s(wfa_s_323), 
       .cout(wfa_cout_323));   // mult.v(3090)
    and (wand_941, a[29], b[13]) ;   // mult.v(3091)
    and (wand_972, a[30], b[12]) ;   // mult.v(3092)
    and (wand_1003, a[31], b[11]) ;   // mult.v(3093)
    fa fa_324 (.a(wand_941), .b(wand_972), .cin(wand_1003), .s(wfa_s_324), 
       .cout(wfa_cout_324));   // mult.v(3094)
    fa fa_325 (.a(wfa_cout_158), .b(wfa_cout_159), .cin(wfa_cout_160), 
       .s(wfa_s_325), .cout(wfa_cout_325));   // mult.v(3095)
    fa fa_326 (.a(wfa_cout_161), .b(wfa_s_162), .cin(wfa_s_163), .s(wfa_s_326), 
       .cout(wfa_cout_326));   // mult.v(3096)
    and (wand_601, a[18], b[25]) ;   // mult.v(3097)
    and (wand_632, a[19], b[24]) ;   // mult.v(3098)
    and (wand_663, a[20], b[23]) ;   // mult.v(3099)
    fa fa_327 (.a(wand_601), .b(wand_632), .cin(wand_663), .s(wfa_s_327), 
       .cout(wfa_cout_327));   // mult.v(3100)
    and (wand_694, a[21], b[22]) ;   // mult.v(3101)
    and (wand_725, a[22], b[21]) ;   // mult.v(3102)
    and (wand_756, a[23], b[20]) ;   // mult.v(3103)
    fa fa_328 (.a(wand_694), .b(wand_725), .cin(wand_756), .s(wfa_s_328), 
       .cout(wfa_cout_328));   // mult.v(3104)
    and (wand_787, a[24], b[19]) ;   // mult.v(3105)
    and (wand_818, a[25], b[18]) ;   // mult.v(3106)
    and (wand_849, a[26], b[17]) ;   // mult.v(3107)
    fa fa_329 (.a(wand_787), .b(wand_818), .cin(wand_849), .s(wfa_s_329), 
       .cout(wfa_cout_329));   // mult.v(3108)
    and (wand_880, a[27], b[16]) ;   // mult.v(3109)
    and (wand_911, a[28], b[15]) ;   // mult.v(3110)
    and (wand_942, a[29], b[14]) ;   // mult.v(3111)
    fa fa_330 (.a(wand_880), .b(wand_911), .cin(wand_942), .s(wfa_s_330), 
       .cout(wfa_cout_330));   // mult.v(3112)
    and (wand_973, a[30], b[13]) ;   // mult.v(3113)
    and (wand_1004, a[31], b[12]) ;   // mult.v(3114)
    fa fa_331 (.a(wand_973), .b(wand_1004), .cin(wfa_cout_162), .s(wfa_s_331), 
       .cout(wfa_cout_331));   // mult.v(3115)
    fa fa_332 (.a(wfa_cout_163), .b(wfa_cout_164), .cin(wfa_s_165), .s(wfa_s_332), 
       .cout(wfa_cout_332));   // mult.v(3116)
    and (wand_540, a[16], b[28]) ;   // mult.v(3117)
    and (wand_571, a[17], b[27]) ;   // mult.v(3118)
    and (wand_602, a[18], b[26]) ;   // mult.v(3119)
    fa fa_333 (.a(wand_540), .b(wand_571), .cin(wand_602), .s(wfa_s_333), 
       .cout(wfa_cout_333));   // mult.v(3120)
    and (wand_633, a[19], b[25]) ;   // mult.v(3121)
    and (wand_664, a[20], b[24]) ;   // mult.v(3122)
    and (wand_695, a[21], b[23]) ;   // mult.v(3123)
    fa fa_334 (.a(wand_633), .b(wand_664), .cin(wand_695), .s(wfa_s_334), 
       .cout(wfa_cout_334));   // mult.v(3124)
    and (wand_726, a[22], b[22]) ;   // mult.v(3125)
    and (wand_757, a[23], b[21]) ;   // mult.v(3126)
    and (wand_788, a[24], b[20]) ;   // mult.v(3127)
    fa fa_335 (.a(wand_726), .b(wand_757), .cin(wand_788), .s(wfa_s_335), 
       .cout(wfa_cout_335));   // mult.v(3128)
    and (wand_819, a[25], b[19]) ;   // mult.v(3129)
    and (wand_850, a[26], b[18]) ;   // mult.v(3130)
    and (wand_881, a[27], b[17]) ;   // mult.v(3131)
    fa fa_336 (.a(wand_819), .b(wand_850), .cin(wand_881), .s(wfa_s_336), 
       .cout(wfa_cout_336));   // mult.v(3132)
    and (wand_912, a[28], b[16]) ;   // mult.v(3133)
    and (wand_943, a[29], b[15]) ;   // mult.v(3134)
    and (wand_974, a[30], b[14]) ;   // mult.v(3135)
    fa fa_337 (.a(wand_912), .b(wand_943), .cin(wand_974), .s(wfa_s_337), 
       .cout(wfa_cout_337));   // mult.v(3136)
    and (wand_1005, a[31], b[13]) ;   // mult.v(3137)
    fa fa_338 (.a(wand_1005), .b(wfa_cout_165), .cin(wfa_cout_166), .s(wfa_s_338), 
       .cout(wfa_cout_338));   // mult.v(3138)
    and (wand_479, a[14], b[31]) ;   // mult.v(3139)
    and (wand_510, a[15], b[30]) ;   // mult.v(3140)
    and (wand_541, a[16], b[29]) ;   // mult.v(3141)
    fa fa_339 (.a(wand_479), .b(wand_510), .cin(wand_541), .s(wfa_s_339), 
       .cout(wfa_cout_339));   // mult.v(3142)
    and (wand_572, a[17], b[28]) ;   // mult.v(3143)
    and (wand_603, a[18], b[27]) ;   // mult.v(3144)
    and (wand_634, a[19], b[26]) ;   // mult.v(3145)
    fa fa_340 (.a(wand_572), .b(wand_603), .cin(wand_634), .s(wfa_s_340), 
       .cout(wfa_cout_340));   // mult.v(3146)
    and (wand_665, a[20], b[25]) ;   // mult.v(3147)
    and (wand_696, a[21], b[24]) ;   // mult.v(3148)
    and (wand_727, a[22], b[23]) ;   // mult.v(3149)
    fa fa_341 (.a(wand_665), .b(wand_696), .cin(wand_727), .s(wfa_s_341), 
       .cout(wfa_cout_341));   // mult.v(3150)
    and (wand_758, a[23], b[22]) ;   // mult.v(3151)
    and (wand_789, a[24], b[21]) ;   // mult.v(3152)
    and (wand_820, a[25], b[20]) ;   // mult.v(3153)
    fa fa_342 (.a(wand_758), .b(wand_789), .cin(wand_820), .s(wfa_s_342), 
       .cout(wfa_cout_342));   // mult.v(3154)
    and (wand_851, a[26], b[19]) ;   // mult.v(3155)
    and (wand_882, a[27], b[18]) ;   // mult.v(3156)
    and (wand_913, a[28], b[17]) ;   // mult.v(3157)
    fa fa_343 (.a(wand_851), .b(wand_882), .cin(wand_913), .s(wfa_s_343), 
       .cout(wfa_cout_343));   // mult.v(3158)
    and (wand_944, a[29], b[16]) ;   // mult.v(3159)
    and (wand_975, a[30], b[15]) ;   // mult.v(3160)
    and (wand_1006, a[31], b[14]) ;   // mult.v(3161)
    fa fa_344 (.a(wand_944), .b(wand_975), .cin(wand_1006), .s(wfa_s_344), 
       .cout(wfa_cout_344));   // mult.v(3162)
    and (wand_511, a[15], b[31]) ;   // mult.v(3163)
    and (wand_542, a[16], b[30]) ;   // mult.v(3164)
    and (wand_573, a[17], b[29]) ;   // mult.v(3165)
    fa fa_345 (.a(wand_511), .b(wand_542), .cin(wand_573), .s(wfa_s_345), 
       .cout(wfa_cout_345));   // mult.v(3166)
    and (wand_604, a[18], b[28]) ;   // mult.v(3167)
    and (wand_635, a[19], b[27]) ;   // mult.v(3168)
    and (wand_666, a[20], b[26]) ;   // mult.v(3169)
    fa fa_346 (.a(wand_604), .b(wand_635), .cin(wand_666), .s(wfa_s_346), 
       .cout(wfa_cout_346));   // mult.v(3170)
    and (wand_697, a[21], b[25]) ;   // mult.v(3171)
    and (wand_728, a[22], b[24]) ;   // mult.v(3172)
    and (wand_759, a[23], b[23]) ;   // mult.v(3173)
    fa fa_347 (.a(wand_697), .b(wand_728), .cin(wand_759), .s(wfa_s_347), 
       .cout(wfa_cout_347));   // mult.v(3174)
    and (wand_790, a[24], b[22]) ;   // mult.v(3175)
    and (wand_821, a[25], b[21]) ;   // mult.v(3176)
    and (wand_852, a[26], b[20]) ;   // mult.v(3177)
    fa fa_348 (.a(wand_790), .b(wand_821), .cin(wand_852), .s(wfa_s_348), 
       .cout(wfa_cout_348));   // mult.v(3178)
    and (wand_883, a[27], b[19]) ;   // mult.v(3179)
    and (wand_914, a[28], b[18]) ;   // mult.v(3180)
    and (wand_945, a[29], b[17]) ;   // mult.v(3181)
    fa fa_349 (.a(wand_883), .b(wand_914), .cin(wand_945), .s(wfa_s_349), 
       .cout(wfa_cout_349));   // mult.v(3182)
    and (wand_543, a[16], b[31]) ;   // mult.v(3183)
    and (wand_574, a[17], b[30]) ;   // mult.v(3184)
    and (wand_605, a[18], b[29]) ;   // mult.v(3185)
    fa fa_350 (.a(wand_543), .b(wand_574), .cin(wand_605), .s(wfa_s_350), 
       .cout(wfa_cout_350));   // mult.v(3186)
    and (wand_636, a[19], b[28]) ;   // mult.v(3187)
    and (wand_667, a[20], b[27]) ;   // mult.v(3188)
    and (wand_698, a[21], b[26]) ;   // mult.v(3189)
    fa fa_351 (.a(wand_636), .b(wand_667), .cin(wand_698), .s(wfa_s_351), 
       .cout(wfa_cout_351));   // mult.v(3190)
    and (wand_729, a[22], b[25]) ;   // mult.v(3191)
    and (wand_760, a[23], b[24]) ;   // mult.v(3192)
    and (wand_791, a[24], b[23]) ;   // mult.v(3193)
    fa fa_352 (.a(wand_729), .b(wand_760), .cin(wand_791), .s(wfa_s_352), 
       .cout(wfa_cout_352));   // mult.v(3194)
    and (wand_822, a[25], b[22]) ;   // mult.v(3195)
    and (wand_853, a[26], b[21]) ;   // mult.v(3196)
    and (wand_884, a[27], b[20]) ;   // mult.v(3197)
    fa fa_353 (.a(wand_822), .b(wand_853), .cin(wand_884), .s(wfa_s_353), 
       .cout(wfa_cout_353));   // mult.v(3198)
    and (wand_575, a[17], b[31]) ;   // mult.v(3199)
    and (wand_606, a[18], b[30]) ;   // mult.v(3200)
    and (wand_637, a[19], b[29]) ;   // mult.v(3201)
    fa fa_354 (.a(wand_575), .b(wand_606), .cin(wand_637), .s(wfa_s_354), 
       .cout(wfa_cout_354));   // mult.v(3202)
    and (wand_668, a[20], b[28]) ;   // mult.v(3203)
    and (wand_699, a[21], b[27]) ;   // mult.v(3204)
    and (wand_730, a[22], b[26]) ;   // mult.v(3205)
    fa fa_355 (.a(wand_668), .b(wand_699), .cin(wand_730), .s(wfa_s_355), 
       .cout(wfa_cout_355));   // mult.v(3206)
    and (wand_761, a[23], b[25]) ;   // mult.v(3207)
    and (wand_792, a[24], b[24]) ;   // mult.v(3208)
    and (wand_823, a[25], b[23]) ;   // mult.v(3209)
    fa fa_356 (.a(wand_761), .b(wand_792), .cin(wand_823), .s(wfa_s_356), 
       .cout(wfa_cout_356));   // mult.v(3210)
    and (wand_607, a[18], b[31]) ;   // mult.v(3211)
    and (wand_638, a[19], b[30]) ;   // mult.v(3212)
    and (wand_669, a[20], b[29]) ;   // mult.v(3213)
    fa fa_357 (.a(wand_607), .b(wand_638), .cin(wand_669), .s(wfa_s_357), 
       .cout(wfa_cout_357));   // mult.v(3214)
    and (wand_700, a[21], b[28]) ;   // mult.v(3215)
    and (wand_731, a[22], b[27]) ;   // mult.v(3216)
    and (wand_762, a[23], b[26]) ;   // mult.v(3217)
    fa fa_358 (.a(wand_700), .b(wand_731), .cin(wand_762), .s(wfa_s_358), 
       .cout(wfa_cout_358));   // mult.v(3218)
    and (wand_639, a[19], b[31]) ;   // mult.v(3219)
    and (wand_670, a[20], b[30]) ;   // mult.v(3220)
    and (wand_701, a[21], b[29]) ;   // mult.v(3221)
    fa fa_359 (.a(wand_639), .b(wand_670), .cin(wand_701), .s(wfa_s_359), 
       .cout(wfa_cout_359));   // mult.v(3222)
    and (wand_9, a[0], b[9]) ;   // mult.v(3223)
    and (wand_40, a[1], b[8]) ;   // mult.v(3224)
    ha ha_20 (.a(wand_9), .b(wand_40), .s(wha_s_20), .c(wha_c_20));   // mult.v(3225)
    and (wand_10, a[0], b[10]) ;   // mult.v(3226)
    and (wand_41, a[1], b[9]) ;   // mult.v(3227)
    and (wand_72, a[2], b[8]) ;   // mult.v(3228)
    fa fa_360 (.a(wand_10), .b(wand_41), .cin(wand_72), .s(wfa_s_360), 
       .cout(wfa_cout_360));   // mult.v(3229)
    and (wand_103, a[3], b[7]) ;   // mult.v(3230)
    and (wand_134, a[4], b[6]) ;   // mult.v(3231)
    ha ha_21 (.a(wand_103), .b(wand_134), .s(wha_s_21), .c(wha_c_21));   // mult.v(3232)
    and (wand_11, a[0], b[11]) ;   // mult.v(3233)
    and (wand_42, a[1], b[10]) ;   // mult.v(3234)
    and (wand_73, a[2], b[9]) ;   // mult.v(3235)
    fa fa_361 (.a(wand_11), .b(wand_42), .cin(wand_73), .s(wfa_s_361), 
       .cout(wfa_cout_361));   // mult.v(3236)
    and (wand_104, a[3], b[8]) ;   // mult.v(3237)
    and (wand_135, a[4], b[7]) ;   // mult.v(3238)
    and (wand_166, a[5], b[6]) ;   // mult.v(3239)
    fa fa_362 (.a(wand_104), .b(wand_135), .cin(wand_166), .s(wfa_s_362), 
       .cout(wfa_cout_362));   // mult.v(3240)
    and (wand_197, a[6], b[5]) ;   // mult.v(3241)
    and (wand_228, a[7], b[4]) ;   // mult.v(3242)
    ha ha_22 (.a(wand_197), .b(wand_228), .s(wha_s_22), .c(wha_c_22));   // mult.v(3243)
    and (wand_12, a[0], b[12]) ;   // mult.v(3244)
    and (wand_43, a[1], b[11]) ;   // mult.v(3245)
    and (wand_74, a[2], b[10]) ;   // mult.v(3246)
    fa fa_363 (.a(wand_12), .b(wand_43), .cin(wand_74), .s(wfa_s_363), 
       .cout(wfa_cout_363));   // mult.v(3247)
    and (wand_105, a[3], b[9]) ;   // mult.v(3248)
    and (wand_136, a[4], b[8]) ;   // mult.v(3249)
    and (wand_167, a[5], b[7]) ;   // mult.v(3250)
    fa fa_364 (.a(wand_105), .b(wand_136), .cin(wand_167), .s(wfa_s_364), 
       .cout(wfa_cout_364));   // mult.v(3251)
    and (wand_198, a[6], b[6]) ;   // mult.v(3252)
    and (wand_229, a[7], b[5]) ;   // mult.v(3253)
    and (wand_260, a[8], b[4]) ;   // mult.v(3254)
    fa fa_365 (.a(wand_198), .b(wand_229), .cin(wand_260), .s(wfa_s_365), 
       .cout(wfa_cout_365));   // mult.v(3255)
    and (wand_291, a[9], b[3]) ;   // mult.v(3256)
    and (wand_322, a[10], b[2]) ;   // mult.v(3257)
    ha ha_23 (.a(wand_291), .b(wand_322), .s(wha_s_23), .c(wha_c_23));   // mult.v(3258)
    and (wand_75, a[2], b[11]) ;   // mult.v(3259)
    and (wand_106, a[3], b[10]) ;   // mult.v(3260)
    and (wand_137, a[4], b[9]) ;   // mult.v(3261)
    fa fa_366 (.a(wand_75), .b(wand_106), .cin(wand_137), .s(wfa_s_366), 
       .cout(wfa_cout_366));   // mult.v(3262)
    and (wand_168, a[5], b[8]) ;   // mult.v(3263)
    and (wand_199, a[6], b[7]) ;   // mult.v(3264)
    and (wand_230, a[7], b[6]) ;   // mult.v(3265)
    fa fa_367 (.a(wand_168), .b(wand_199), .cin(wand_230), .s(wfa_s_367), 
       .cout(wfa_cout_367));   // mult.v(3266)
    and (wand_261, a[8], b[5]) ;   // mult.v(3267)
    and (wand_292, a[9], b[4]) ;   // mult.v(3268)
    and (wand_323, a[10], b[3]) ;   // mult.v(3269)
    fa fa_368 (.a(wand_261), .b(wand_292), .cin(wand_323), .s(wfa_s_368), 
       .cout(wfa_cout_368));   // mult.v(3270)
    and (wand_354, a[11], b[2]) ;   // mult.v(3271)
    and (wand_385, a[12], b[1]) ;   // mult.v(3272)
    and (wand_416, a[13], b[0]) ;   // mult.v(3273)
    fa fa_369 (.a(wand_354), .b(wand_385), .cin(wand_416), .s(wfa_s_369), 
       .cout(wfa_cout_369));   // mult.v(3274)
    and (wand_169, a[5], b[9]) ;   // mult.v(3275)
    and (wand_200, a[6], b[8]) ;   // mult.v(3276)
    and (wand_231, a[7], b[7]) ;   // mult.v(3277)
    fa fa_370 (.a(wand_169), .b(wand_200), .cin(wand_231), .s(wfa_s_370), 
       .cout(wfa_cout_370));   // mult.v(3278)
    and (wand_262, a[8], b[6]) ;   // mult.v(3279)
    and (wand_293, a[9], b[5]) ;   // mult.v(3280)
    and (wand_324, a[10], b[4]) ;   // mult.v(3281)
    fa fa_371 (.a(wand_262), .b(wand_293), .cin(wand_324), .s(wfa_s_371), 
       .cout(wfa_cout_371));   // mult.v(3282)
    and (wand_355, a[11], b[3]) ;   // mult.v(3283)
    and (wand_386, a[12], b[2]) ;   // mult.v(3284)
    and (wand_417, a[13], b[1]) ;   // mult.v(3285)
    fa fa_372 (.a(wand_355), .b(wand_386), .cin(wand_417), .s(wfa_s_372), 
       .cout(wfa_cout_372));   // mult.v(3286)
    and (wand_448, a[14], b[0]) ;   // mult.v(3287)
    fa fa_373 (.a(wand_448), .b(wha_c_14), .cin(wfa_s_168), .s(wfa_s_373), 
       .cout(wfa_cout_373));   // mult.v(3288)
    and (wand_263, a[8], b[7]) ;   // mult.v(3289)
    and (wand_294, a[9], b[6]) ;   // mult.v(3290)
    and (wand_325, a[10], b[5]) ;   // mult.v(3291)
    fa fa_374 (.a(wand_263), .b(wand_294), .cin(wand_325), .s(wfa_s_374), 
       .cout(wfa_cout_374));   // mult.v(3292)
    and (wand_356, a[11], b[4]) ;   // mult.v(3293)
    and (wand_387, a[12], b[3]) ;   // mult.v(3294)
    and (wand_418, a[13], b[2]) ;   // mult.v(3295)
    fa fa_375 (.a(wand_356), .b(wand_387), .cin(wand_418), .s(wfa_s_375), 
       .cout(wfa_cout_375));   // mult.v(3296)
    and (wand_449, a[14], b[1]) ;   // mult.v(3297)
    and (wand_480, a[15], b[0]) ;   // mult.v(3298)
    fa fa_376 (.a(wand_449), .b(wand_480), .cin(wfa_cout_168), .s(wfa_s_376), 
       .cout(wfa_cout_376));   // mult.v(3299)
    fa fa_377 (.a(wha_c_15), .b(wfa_s_169), .cin(wfa_s_170), .s(wfa_s_377), 
       .cout(wfa_cout_377));   // mult.v(3300)
    and (wand_357, a[11], b[5]) ;   // mult.v(3301)
    and (wand_388, a[12], b[4]) ;   // mult.v(3302)
    and (wand_419, a[13], b[3]) ;   // mult.v(3303)
    fa fa_378 (.a(wand_357), .b(wand_388), .cin(wand_419), .s(wfa_s_378), 
       .cout(wfa_cout_378));   // mult.v(3304)
    and (wand_450, a[14], b[2]) ;   // mult.v(3305)
    and (wand_481, a[15], b[1]) ;   // mult.v(3306)
    and (wand_512, a[16], b[0]) ;   // mult.v(3307)
    fa fa_379 (.a(wand_450), .b(wand_481), .cin(wand_512), .s(wfa_s_379), 
       .cout(wfa_cout_379));   // mult.v(3308)
    fa fa_380 (.a(wfa_cout_169), .b(wfa_cout_170), .cin(wha_c_16), .s(wfa_s_380), 
       .cout(wfa_cout_380));   // mult.v(3309)
    fa fa_381 (.a(wfa_s_171), .b(wfa_s_172), .cin(wfa_s_173), .s(wfa_s_381), 
       .cout(wfa_cout_381));   // mult.v(3310)
    and (wand_451, a[14], b[3]) ;   // mult.v(3311)
    and (wand_482, a[15], b[2]) ;   // mult.v(3312)
    and (wand_513, a[16], b[1]) ;   // mult.v(3313)
    fa fa_382 (.a(wand_451), .b(wand_482), .cin(wand_513), .s(wfa_s_382), 
       .cout(wfa_cout_382));   // mult.v(3314)
    and (wand_544, a[17], b[0]) ;   // mult.v(3315)
    fa fa_383 (.a(wand_544), .b(wfa_cout_171), .cin(wfa_cout_172), .s(wfa_s_383), 
       .cout(wfa_cout_383));   // mult.v(3316)
    fa fa_384 (.a(wfa_cout_173), .b(wha_c_17), .cin(wfa_s_174), .s(wfa_s_384), 
       .cout(wfa_cout_384));   // mult.v(3317)
    fa fa_385 (.a(wfa_s_175), .b(wfa_s_176), .cin(wfa_s_177), .s(wfa_s_385), 
       .cout(wfa_cout_385));   // mult.v(3318)
    and (wand_545, a[17], b[1]) ;   // mult.v(3319)
    and (wand_576, a[18], b[0]) ;   // mult.v(3320)
    fa fa_386 (.a(wand_545), .b(wand_576), .cin(wfa_cout_174), .s(wfa_s_386), 
       .cout(wfa_cout_386));   // mult.v(3321)
    fa fa_387 (.a(wfa_cout_175), .b(wfa_cout_176), .cin(wfa_cout_177), 
       .s(wfa_s_387), .cout(wfa_cout_387));   // mult.v(3322)
    fa fa_388 (.a(wha_c_18), .b(wfa_s_178), .cin(wfa_s_179), .s(wfa_s_388), 
       .cout(wfa_cout_388));   // mult.v(3323)
    fa fa_389 (.a(wfa_s_180), .b(wfa_s_181), .cin(wfa_s_182), .s(wfa_s_389), 
       .cout(wfa_cout_389));   // mult.v(3324)
    fa fa_390 (.a(wha_s_5), .b(wfa_cout_178), .cin(wfa_cout_179), .s(wfa_s_390), 
       .cout(wfa_cout_390));   // mult.v(3325)
    fa fa_391 (.a(wfa_cout_180), .b(wfa_cout_181), .cin(wfa_cout_182), 
       .s(wfa_s_391), .cout(wfa_cout_391));   // mult.v(3326)
    fa fa_392 (.a(wha_c_19), .b(wfa_s_183), .cin(wfa_s_184), .s(wfa_s_392), 
       .cout(wfa_cout_392));   // mult.v(3327)
    fa fa_393 (.a(wfa_s_185), .b(wfa_s_186), .cin(wfa_s_187), .s(wfa_s_393), 
       .cout(wfa_cout_393));   // mult.v(3328)
    fa fa_394 (.a(wha_s_6), .b(wfa_cout_183), .cin(wfa_cout_184), .s(wfa_s_394), 
       .cout(wfa_cout_394));   // mult.v(3329)
    fa fa_395 (.a(wfa_cout_185), .b(wfa_cout_186), .cin(wfa_cout_187), 
       .s(wfa_s_395), .cout(wfa_cout_395));   // mult.v(3330)
    fa fa_396 (.a(wfa_cout_188), .b(wfa_s_189), .cin(wfa_s_190), .s(wfa_s_396), 
       .cout(wfa_cout_396));   // mult.v(3331)
    fa fa_397 (.a(wfa_s_191), .b(wfa_s_192), .cin(wfa_s_193), .s(wfa_s_397), 
       .cout(wfa_cout_397));   // mult.v(3332)
    fa fa_398 (.a(wha_s_7), .b(wfa_cout_189), .cin(wfa_cout_190), .s(wfa_s_398), 
       .cout(wfa_cout_398));   // mult.v(3333)
    fa fa_399 (.a(wfa_cout_191), .b(wfa_cout_192), .cin(wfa_cout_193), 
       .s(wfa_s_399), .cout(wfa_cout_399));   // mult.v(3334)
    fa fa_400 (.a(wfa_cout_194), .b(wfa_s_195), .cin(wfa_s_196), .s(wfa_s_400), 
       .cout(wfa_cout_400));   // mult.v(3335)
    fa fa_401 (.a(wfa_s_197), .b(wfa_s_198), .cin(wfa_s_199), .s(wfa_s_401), 
       .cout(wfa_cout_401));   // mult.v(3336)
    fa fa_402 (.a(wha_s_8), .b(wfa_cout_195), .cin(wfa_cout_196), .s(wfa_s_402), 
       .cout(wfa_cout_402));   // mult.v(3337)
    fa fa_403 (.a(wfa_cout_197), .b(wfa_cout_198), .cin(wfa_cout_199), 
       .s(wfa_s_403), .cout(wfa_cout_403));   // mult.v(3338)
    fa fa_404 (.a(wfa_cout_200), .b(wfa_s_201), .cin(wfa_s_202), .s(wfa_s_404), 
       .cout(wfa_cout_404));   // mult.v(3339)
    fa fa_405 (.a(wfa_s_203), .b(wfa_s_204), .cin(wfa_s_205), .s(wfa_s_405), 
       .cout(wfa_cout_405));   // mult.v(3340)
    fa fa_406 (.a(wha_s_9), .b(wfa_cout_201), .cin(wfa_cout_202), .s(wfa_s_406), 
       .cout(wfa_cout_406));   // mult.v(3341)
    fa fa_407 (.a(wfa_cout_203), .b(wfa_cout_204), .cin(wfa_cout_205), 
       .s(wfa_s_407), .cout(wfa_cout_407));   // mult.v(3342)
    fa fa_408 (.a(wfa_cout_206), .b(wfa_s_207), .cin(wfa_s_208), .s(wfa_s_408), 
       .cout(wfa_cout_408));   // mult.v(3343)
    fa fa_409 (.a(wfa_s_209), .b(wfa_s_210), .cin(wfa_s_211), .s(wfa_s_409), 
       .cout(wfa_cout_409));   // mult.v(3344)
    fa fa_410 (.a(wha_s_10), .b(wfa_cout_207), .cin(wfa_cout_208), .s(wfa_s_410), 
       .cout(wfa_cout_410));   // mult.v(3345)
    fa fa_411 (.a(wfa_cout_209), .b(wfa_cout_210), .cin(wfa_cout_211), 
       .s(wfa_s_411), .cout(wfa_cout_411));   // mult.v(3346)
    fa fa_412 (.a(wfa_cout_212), .b(wfa_s_213), .cin(wfa_s_214), .s(wfa_s_412), 
       .cout(wfa_cout_412));   // mult.v(3347)
    fa fa_413 (.a(wfa_s_215), .b(wfa_s_216), .cin(wfa_s_217), .s(wfa_s_413), 
       .cout(wfa_cout_413));   // mult.v(3348)
    fa fa_414 (.a(wha_s_11), .b(wfa_cout_213), .cin(wfa_cout_214), .s(wfa_s_414), 
       .cout(wfa_cout_414));   // mult.v(3349)
    fa fa_415 (.a(wfa_cout_215), .b(wfa_cout_216), .cin(wfa_cout_217), 
       .s(wfa_s_415), .cout(wfa_cout_415));   // mult.v(3350)
    fa fa_416 (.a(wfa_cout_218), .b(wfa_s_219), .cin(wfa_s_220), .s(wfa_s_416), 
       .cout(wfa_cout_416));   // mult.v(3351)
    fa fa_417 (.a(wfa_s_221), .b(wfa_s_222), .cin(wfa_s_223), .s(wfa_s_417), 
       .cout(wfa_cout_417));   // mult.v(3352)
    fa fa_418 (.a(wha_s_12), .b(wfa_cout_219), .cin(wfa_cout_220), .s(wfa_s_418), 
       .cout(wfa_cout_418));   // mult.v(3353)
    fa fa_419 (.a(wfa_cout_221), .b(wfa_cout_222), .cin(wfa_cout_223), 
       .s(wfa_s_419), .cout(wfa_cout_419));   // mult.v(3354)
    fa fa_420 (.a(wfa_cout_224), .b(wfa_s_225), .cin(wfa_s_226), .s(wfa_s_420), 
       .cout(wfa_cout_420));   // mult.v(3355)
    fa fa_421 (.a(wfa_s_227), .b(wfa_s_228), .cin(wfa_s_229), .s(wfa_s_421), 
       .cout(wfa_cout_421));   // mult.v(3356)
    fa fa_422 (.a(wha_s_13), .b(wfa_cout_225), .cin(wfa_cout_226), .s(wfa_s_422), 
       .cout(wfa_cout_422));   // mult.v(3357)
    fa fa_423 (.a(wfa_cout_227), .b(wfa_cout_228), .cin(wfa_cout_229), 
       .s(wfa_s_423), .cout(wfa_cout_423));   // mult.v(3358)
    fa fa_424 (.a(wfa_cout_230), .b(wfa_s_231), .cin(wfa_s_232), .s(wfa_s_424), 
       .cout(wfa_cout_424));   // mult.v(3359)
    fa fa_425 (.a(wfa_s_233), .b(wfa_s_234), .cin(wfa_s_235), .s(wfa_s_425), 
       .cout(wfa_cout_425));   // mult.v(3360)
    fa fa_426 (.a(wfa_s_59), .b(wfa_cout_231), .cin(wfa_cout_232), .s(wfa_s_426), 
       .cout(wfa_cout_426));   // mult.v(3361)
    fa fa_427 (.a(wfa_cout_233), .b(wfa_cout_234), .cin(wfa_cout_235), 
       .s(wfa_s_427), .cout(wfa_cout_427));   // mult.v(3362)
    fa fa_428 (.a(wfa_cout_236), .b(wfa_s_237), .cin(wfa_s_238), .s(wfa_s_428), 
       .cout(wfa_cout_428));   // mult.v(3363)
    fa fa_429 (.a(wfa_s_239), .b(wfa_s_240), .cin(wfa_s_241), .s(wfa_s_429), 
       .cout(wfa_cout_429));   // mult.v(3364)
    fa fa_430 (.a(wfa_s_68), .b(wfa_cout_237), .cin(wfa_cout_238), .s(wfa_s_430), 
       .cout(wfa_cout_430));   // mult.v(3365)
    fa fa_431 (.a(wfa_cout_239), .b(wfa_cout_240), .cin(wfa_cout_241), 
       .s(wfa_s_431), .cout(wfa_cout_431));   // mult.v(3366)
    fa fa_432 (.a(wfa_cout_242), .b(wfa_s_243), .cin(wfa_s_244), .s(wfa_s_432), 
       .cout(wfa_cout_432));   // mult.v(3367)
    fa fa_433 (.a(wfa_s_245), .b(wfa_s_246), .cin(wfa_s_247), .s(wfa_s_433), 
       .cout(wfa_cout_433));   // mult.v(3368)
    fa fa_434 (.a(wfa_s_77), .b(wfa_cout_243), .cin(wfa_cout_244), .s(wfa_s_434), 
       .cout(wfa_cout_434));   // mult.v(3369)
    fa fa_435 (.a(wfa_cout_245), .b(wfa_cout_246), .cin(wfa_cout_247), 
       .s(wfa_s_435), .cout(wfa_cout_435));   // mult.v(3370)
    fa fa_436 (.a(wfa_cout_248), .b(wfa_s_249), .cin(wfa_s_250), .s(wfa_s_436), 
       .cout(wfa_cout_436));   // mult.v(3371)
    fa fa_437 (.a(wfa_s_251), .b(wfa_s_252), .cin(wfa_s_253), .s(wfa_s_437), 
       .cout(wfa_cout_437));   // mult.v(3372)
    fa fa_438 (.a(wfa_s_86), .b(wfa_cout_249), .cin(wfa_cout_250), .s(wfa_s_438), 
       .cout(wfa_cout_438));   // mult.v(3373)
    fa fa_439 (.a(wfa_cout_251), .b(wfa_cout_252), .cin(wfa_cout_253), 
       .s(wfa_s_439), .cout(wfa_cout_439));   // mult.v(3374)
    fa fa_440 (.a(wfa_cout_254), .b(wfa_s_255), .cin(wfa_s_256), .s(wfa_s_440), 
       .cout(wfa_cout_440));   // mult.v(3375)
    fa fa_441 (.a(wfa_s_257), .b(wfa_s_258), .cin(wfa_s_259), .s(wfa_s_441), 
       .cout(wfa_cout_441));   // mult.v(3376)
    fa fa_442 (.a(wfa_s_95), .b(wfa_cout_255), .cin(wfa_cout_256), .s(wfa_s_442), 
       .cout(wfa_cout_442));   // mult.v(3377)
    fa fa_443 (.a(wfa_cout_257), .b(wfa_cout_258), .cin(wfa_cout_259), 
       .s(wfa_s_443), .cout(wfa_cout_443));   // mult.v(3378)
    fa fa_444 (.a(wfa_cout_260), .b(wfa_s_261), .cin(wfa_s_262), .s(wfa_s_444), 
       .cout(wfa_cout_444));   // mult.v(3379)
    fa fa_445 (.a(wfa_s_263), .b(wfa_s_264), .cin(wfa_s_265), .s(wfa_s_445), 
       .cout(wfa_cout_445));   // mult.v(3380)
    fa fa_446 (.a(wfa_s_104), .b(wfa_cout_261), .cin(wfa_cout_262), .s(wfa_s_446), 
       .cout(wfa_cout_446));   // mult.v(3381)
    fa fa_447 (.a(wfa_cout_263), .b(wfa_cout_264), .cin(wfa_cout_265), 
       .s(wfa_s_447), .cout(wfa_cout_447));   // mult.v(3382)
    fa fa_448 (.a(wfa_cout_266), .b(wfa_s_267), .cin(wfa_s_268), .s(wfa_s_448), 
       .cout(wfa_cout_448));   // mult.v(3383)
    fa fa_449 (.a(wfa_s_269), .b(wfa_s_270), .cin(wfa_s_271), .s(wfa_s_449), 
       .cout(wfa_cout_449));   // mult.v(3384)
    fa fa_450 (.a(wfa_s_113), .b(wfa_cout_267), .cin(wfa_cout_268), .s(wfa_s_450), 
       .cout(wfa_cout_450));   // mult.v(3385)
    fa fa_451 (.a(wfa_cout_269), .b(wfa_cout_270), .cin(wfa_cout_271), 
       .s(wfa_s_451), .cout(wfa_cout_451));   // mult.v(3386)
    fa fa_452 (.a(wfa_cout_272), .b(wfa_s_273), .cin(wfa_s_274), .s(wfa_s_452), 
       .cout(wfa_cout_452));   // mult.v(3387)
    fa fa_453 (.a(wfa_s_275), .b(wfa_s_276), .cin(wfa_s_277), .s(wfa_s_453), 
       .cout(wfa_cout_453));   // mult.v(3388)
    fa fa_454 (.a(wfa_s_122), .b(wfa_cout_273), .cin(wfa_cout_274), .s(wfa_s_454), 
       .cout(wfa_cout_454));   // mult.v(3389)
    fa fa_455 (.a(wfa_cout_275), .b(wfa_cout_276), .cin(wfa_cout_277), 
       .s(wfa_s_455), .cout(wfa_cout_455));   // mult.v(3390)
    fa fa_456 (.a(wfa_cout_278), .b(wfa_s_279), .cin(wfa_s_280), .s(wfa_s_456), 
       .cout(wfa_cout_456));   // mult.v(3391)
    fa fa_457 (.a(wfa_s_281), .b(wfa_s_282), .cin(wfa_s_283), .s(wfa_s_457), 
       .cout(wfa_cout_457));   // mult.v(3392)
    fa fa_458 (.a(wfa_s_131), .b(wfa_cout_279), .cin(wfa_cout_280), .s(wfa_s_458), 
       .cout(wfa_cout_458));   // mult.v(3393)
    fa fa_459 (.a(wfa_cout_281), .b(wfa_cout_282), .cin(wfa_cout_283), 
       .s(wfa_s_459), .cout(wfa_cout_459));   // mult.v(3394)
    fa fa_460 (.a(wfa_cout_284), .b(wfa_s_285), .cin(wfa_s_286), .s(wfa_s_460), 
       .cout(wfa_cout_460));   // mult.v(3395)
    fa fa_461 (.a(wfa_s_287), .b(wfa_s_288), .cin(wfa_s_289), .s(wfa_s_461), 
       .cout(wfa_cout_461));   // mult.v(3396)
    fa fa_462 (.a(wfa_s_139), .b(wfa_cout_285), .cin(wfa_cout_286), .s(wfa_s_462), 
       .cout(wfa_cout_462));   // mult.v(3397)
    fa fa_463 (.a(wfa_cout_287), .b(wfa_cout_288), .cin(wfa_cout_289), 
       .s(wfa_s_463), .cout(wfa_cout_463));   // mult.v(3398)
    fa fa_464 (.a(wfa_cout_290), .b(wfa_s_291), .cin(wfa_s_292), .s(wfa_s_464), 
       .cout(wfa_cout_464));   // mult.v(3399)
    fa fa_465 (.a(wfa_s_293), .b(wfa_s_294), .cin(wfa_s_295), .s(wfa_s_465), 
       .cout(wfa_cout_465));   // mult.v(3400)
    fa fa_466 (.a(wfa_s_146), .b(wfa_cout_291), .cin(wfa_cout_292), .s(wfa_s_466), 
       .cout(wfa_cout_466));   // mult.v(3401)
    fa fa_467 (.a(wfa_cout_293), .b(wfa_cout_294), .cin(wfa_cout_295), 
       .s(wfa_s_467), .cout(wfa_cout_467));   // mult.v(3402)
    fa fa_468 (.a(wfa_cout_296), .b(wfa_s_297), .cin(wfa_s_298), .s(wfa_s_468), 
       .cout(wfa_cout_468));   // mult.v(3403)
    fa fa_469 (.a(wfa_s_299), .b(wfa_s_300), .cin(wfa_s_301), .s(wfa_s_469), 
       .cout(wfa_cout_469));   // mult.v(3404)
    fa fa_470 (.a(wfa_s_152), .b(wfa_cout_297), .cin(wfa_cout_298), .s(wfa_s_470), 
       .cout(wfa_cout_470));   // mult.v(3405)
    fa fa_471 (.a(wfa_cout_299), .b(wfa_cout_300), .cin(wfa_cout_301), 
       .s(wfa_s_471), .cout(wfa_cout_471));   // mult.v(3406)
    fa fa_472 (.a(wfa_cout_302), .b(wfa_s_303), .cin(wfa_s_304), .s(wfa_s_472), 
       .cout(wfa_cout_472));   // mult.v(3407)
    fa fa_473 (.a(wfa_s_305), .b(wfa_s_306), .cin(wfa_s_307), .s(wfa_s_473), 
       .cout(wfa_cout_473));   // mult.v(3408)
    fa fa_474 (.a(wfa_s_157), .b(wfa_cout_303), .cin(wfa_cout_304), .s(wfa_s_474), 
       .cout(wfa_cout_474));   // mult.v(3409)
    fa fa_475 (.a(wfa_cout_305), .b(wfa_cout_306), .cin(wfa_cout_307), 
       .s(wfa_s_475), .cout(wfa_cout_475));   // mult.v(3410)
    fa fa_476 (.a(wfa_cout_308), .b(wfa_s_309), .cin(wfa_s_310), .s(wfa_s_476), 
       .cout(wfa_cout_476));   // mult.v(3411)
    fa fa_477 (.a(wfa_s_311), .b(wfa_s_312), .cin(wfa_s_313), .s(wfa_s_477), 
       .cout(wfa_cout_477));   // mult.v(3412)
    fa fa_478 (.a(wfa_s_161), .b(wfa_cout_309), .cin(wfa_cout_310), .s(wfa_s_478), 
       .cout(wfa_cout_478));   // mult.v(3413)
    fa fa_479 (.a(wfa_cout_311), .b(wfa_cout_312), .cin(wfa_cout_313), 
       .s(wfa_s_479), .cout(wfa_cout_479));   // mult.v(3414)
    fa fa_480 (.a(wfa_cout_314), .b(wfa_s_315), .cin(wfa_s_316), .s(wfa_s_480), 
       .cout(wfa_cout_480));   // mult.v(3415)
    fa fa_481 (.a(wfa_s_317), .b(wfa_s_318), .cin(wfa_s_319), .s(wfa_s_481), 
       .cout(wfa_cout_481));   // mult.v(3416)
    fa fa_482 (.a(wfa_s_164), .b(wfa_cout_315), .cin(wfa_cout_316), .s(wfa_s_482), 
       .cout(wfa_cout_482));   // mult.v(3417)
    fa fa_483 (.a(wfa_cout_317), .b(wfa_cout_318), .cin(wfa_cout_319), 
       .s(wfa_s_483), .cout(wfa_cout_483));   // mult.v(3418)
    fa fa_484 (.a(wfa_cout_320), .b(wfa_s_321), .cin(wfa_s_322), .s(wfa_s_484), 
       .cout(wfa_cout_484));   // mult.v(3419)
    fa fa_485 (.a(wfa_s_323), .b(wfa_s_324), .cin(wfa_s_325), .s(wfa_s_485), 
       .cout(wfa_cout_485));   // mult.v(3420)
    fa fa_486 (.a(wfa_s_166), .b(wfa_cout_321), .cin(wfa_cout_322), .s(wfa_s_486), 
       .cout(wfa_cout_486));   // mult.v(3421)
    fa fa_487 (.a(wfa_cout_323), .b(wfa_cout_324), .cin(wfa_cout_325), 
       .s(wfa_s_487), .cout(wfa_cout_487));   // mult.v(3422)
    fa fa_488 (.a(wfa_cout_326), .b(wfa_s_327), .cin(wfa_s_328), .s(wfa_s_488), 
       .cout(wfa_cout_488));   // mult.v(3423)
    fa fa_489 (.a(wfa_s_329), .b(wfa_s_330), .cin(wfa_s_331), .s(wfa_s_489), 
       .cout(wfa_cout_489));   // mult.v(3424)
    fa fa_490 (.a(wfa_s_167), .b(wfa_cout_327), .cin(wfa_cout_328), .s(wfa_s_490), 
       .cout(wfa_cout_490));   // mult.v(3425)
    fa fa_491 (.a(wfa_cout_329), .b(wfa_cout_330), .cin(wfa_cout_331), 
       .s(wfa_s_491), .cout(wfa_cout_491));   // mult.v(3426)
    fa fa_492 (.a(wfa_cout_332), .b(wfa_s_333), .cin(wfa_s_334), .s(wfa_s_492), 
       .cout(wfa_cout_492));   // mult.v(3427)
    fa fa_493 (.a(wfa_s_335), .b(wfa_s_336), .cin(wfa_s_337), .s(wfa_s_493), 
       .cout(wfa_cout_493));   // mult.v(3428)
    fa fa_494 (.a(wfa_cout_167), .b(wfa_cout_333), .cin(wfa_cout_334), 
       .s(wfa_s_494), .cout(wfa_cout_494));   // mult.v(3429)
    fa fa_495 (.a(wfa_cout_335), .b(wfa_cout_336), .cin(wfa_cout_337), 
       .s(wfa_s_495), .cout(wfa_cout_495));   // mult.v(3430)
    fa fa_496 (.a(wfa_cout_338), .b(wfa_s_339), .cin(wfa_s_340), .s(wfa_s_496), 
       .cout(wfa_cout_496));   // mult.v(3431)
    fa fa_497 (.a(wfa_s_341), .b(wfa_s_342), .cin(wfa_s_343), .s(wfa_s_497), 
       .cout(wfa_cout_497));   // mult.v(3432)
    and (wand_976, a[30], b[16]) ;   // mult.v(3433)
    and (wand_1007, a[31], b[15]) ;   // mult.v(3434)
    fa fa_498 (.a(wand_976), .b(wand_1007), .cin(wfa_cout_339), .s(wfa_s_498), 
       .cout(wfa_cout_498));   // mult.v(3435)
    fa fa_499 (.a(wfa_cout_340), .b(wfa_cout_341), .cin(wfa_cout_342), 
       .s(wfa_s_499), .cout(wfa_cout_499));   // mult.v(3436)
    fa fa_500 (.a(wfa_cout_343), .b(wfa_cout_344), .cin(wfa_s_345), .s(wfa_s_500), 
       .cout(wfa_cout_500));   // mult.v(3437)
    fa fa_501 (.a(wfa_s_346), .b(wfa_s_347), .cin(wfa_s_348), .s(wfa_s_501), 
       .cout(wfa_cout_501));   // mult.v(3438)
    and (wand_915, a[28], b[19]) ;   // mult.v(3439)
    and (wand_946, a[29], b[18]) ;   // mult.v(3440)
    and (wand_977, a[30], b[17]) ;   // mult.v(3441)
    fa fa_502 (.a(wand_915), .b(wand_946), .cin(wand_977), .s(wfa_s_502), 
       .cout(wfa_cout_502));   // mult.v(3442)
    and (wand_1008, a[31], b[16]) ;   // mult.v(3443)
    fa fa_503 (.a(wand_1008), .b(wfa_cout_345), .cin(wfa_cout_346), .s(wfa_s_503), 
       .cout(wfa_cout_503));   // mult.v(3444)
    fa fa_504 (.a(wfa_cout_347), .b(wfa_cout_348), .cin(wfa_cout_349), 
       .s(wfa_s_504), .cout(wfa_cout_504));   // mult.v(3445)
    fa fa_505 (.a(wfa_s_350), .b(wfa_s_351), .cin(wfa_s_352), .s(wfa_s_505), 
       .cout(wfa_cout_505));   // mult.v(3446)
    and (wand_854, a[26], b[22]) ;   // mult.v(3447)
    and (wand_885, a[27], b[21]) ;   // mult.v(3448)
    and (wand_916, a[28], b[20]) ;   // mult.v(3449)
    fa fa_506 (.a(wand_854), .b(wand_885), .cin(wand_916), .s(wfa_s_506), 
       .cout(wfa_cout_506));   // mult.v(3450)
    and (wand_947, a[29], b[19]) ;   // mult.v(3451)
    and (wand_978, a[30], b[18]) ;   // mult.v(3452)
    and (wand_1009, a[31], b[17]) ;   // mult.v(3453)
    fa fa_507 (.a(wand_947), .b(wand_978), .cin(wand_1009), .s(wfa_s_507), 
       .cout(wfa_cout_507));   // mult.v(3454)
    fa fa_508 (.a(wfa_cout_350), .b(wfa_cout_351), .cin(wfa_cout_352), 
       .s(wfa_s_508), .cout(wfa_cout_508));   // mult.v(3455)
    fa fa_509 (.a(wfa_cout_353), .b(wfa_s_354), .cin(wfa_s_355), .s(wfa_s_509), 
       .cout(wfa_cout_509));   // mult.v(3456)
    and (wand_793, a[24], b[25]) ;   // mult.v(3457)
    and (wand_824, a[25], b[24]) ;   // mult.v(3458)
    and (wand_855, a[26], b[23]) ;   // mult.v(3459)
    fa fa_510 (.a(wand_793), .b(wand_824), .cin(wand_855), .s(wfa_s_510), 
       .cout(wfa_cout_510));   // mult.v(3460)
    and (wand_886, a[27], b[22]) ;   // mult.v(3461)
    and (wand_917, a[28], b[21]) ;   // mult.v(3462)
    and (wand_948, a[29], b[20]) ;   // mult.v(3463)
    fa fa_511 (.a(wand_886), .b(wand_917), .cin(wand_948), .s(wfa_s_511), 
       .cout(wfa_cout_511));   // mult.v(3464)
    and (wand_979, a[30], b[19]) ;   // mult.v(3465)
    and (wand_1010, a[31], b[18]) ;   // mult.v(3466)
    fa fa_512 (.a(wand_979), .b(wand_1010), .cin(wfa_cout_354), .s(wfa_s_512), 
       .cout(wfa_cout_512));   // mult.v(3467)
    fa fa_513 (.a(wfa_cout_355), .b(wfa_cout_356), .cin(wfa_s_357), .s(wfa_s_513), 
       .cout(wfa_cout_513));   // mult.v(3468)
    and (wand_732, a[22], b[28]) ;   // mult.v(3469)
    and (wand_763, a[23], b[27]) ;   // mult.v(3470)
    and (wand_794, a[24], b[26]) ;   // mult.v(3471)
    fa fa_514 (.a(wand_732), .b(wand_763), .cin(wand_794), .s(wfa_s_514), 
       .cout(wfa_cout_514));   // mult.v(3472)
    and (wand_825, a[25], b[25]) ;   // mult.v(3473)
    and (wand_856, a[26], b[24]) ;   // mult.v(3474)
    and (wand_887, a[27], b[23]) ;   // mult.v(3475)
    fa fa_515 (.a(wand_825), .b(wand_856), .cin(wand_887), .s(wfa_s_515), 
       .cout(wfa_cout_515));   // mult.v(3476)
    and (wand_918, a[28], b[22]) ;   // mult.v(3477)
    and (wand_949, a[29], b[21]) ;   // mult.v(3478)
    and (wand_980, a[30], b[20]) ;   // mult.v(3479)
    fa fa_516 (.a(wand_918), .b(wand_949), .cin(wand_980), .s(wfa_s_516), 
       .cout(wfa_cout_516));   // mult.v(3480)
    and (wand_1011, a[31], b[19]) ;   // mult.v(3481)
    fa fa_517 (.a(wand_1011), .b(wfa_cout_357), .cin(wfa_cout_358), .s(wfa_s_517), 
       .cout(wfa_cout_517));   // mult.v(3482)
    and (wand_671, a[20], b[31]) ;   // mult.v(3483)
    and (wand_702, a[21], b[30]) ;   // mult.v(3484)
    and (wand_733, a[22], b[29]) ;   // mult.v(3485)
    fa fa_518 (.a(wand_671), .b(wand_702), .cin(wand_733), .s(wfa_s_518), 
       .cout(wfa_cout_518));   // mult.v(3486)
    and (wand_764, a[23], b[28]) ;   // mult.v(3487)
    and (wand_795, a[24], b[27]) ;   // mult.v(3488)
    and (wand_826, a[25], b[26]) ;   // mult.v(3489)
    fa fa_519 (.a(wand_764), .b(wand_795), .cin(wand_826), .s(wfa_s_519), 
       .cout(wfa_cout_519));   // mult.v(3490)
    and (wand_857, a[26], b[25]) ;   // mult.v(3491)
    and (wand_888, a[27], b[24]) ;   // mult.v(3492)
    and (wand_919, a[28], b[23]) ;   // mult.v(3493)
    fa fa_520 (.a(wand_857), .b(wand_888), .cin(wand_919), .s(wfa_s_520), 
       .cout(wfa_cout_520));   // mult.v(3494)
    and (wand_950, a[29], b[22]) ;   // mult.v(3495)
    and (wand_981, a[30], b[21]) ;   // mult.v(3496)
    and (wand_1012, a[31], b[20]) ;   // mult.v(3497)
    fa fa_521 (.a(wand_950), .b(wand_981), .cin(wand_1012), .s(wfa_s_521), 
       .cout(wfa_cout_521));   // mult.v(3498)
    and (wand_703, a[21], b[31]) ;   // mult.v(3499)
    and (wand_734, a[22], b[30]) ;   // mult.v(3500)
    and (wand_765, a[23], b[29]) ;   // mult.v(3501)
    fa fa_522 (.a(wand_703), .b(wand_734), .cin(wand_765), .s(wfa_s_522), 
       .cout(wfa_cout_522));   // mult.v(3502)
    and (wand_796, a[24], b[28]) ;   // mult.v(3503)
    and (wand_827, a[25], b[27]) ;   // mult.v(3504)
    and (wand_858, a[26], b[26]) ;   // mult.v(3505)
    fa fa_523 (.a(wand_796), .b(wand_827), .cin(wand_858), .s(wfa_s_523), 
       .cout(wfa_cout_523));   // mult.v(3506)
    and (wand_889, a[27], b[25]) ;   // mult.v(3507)
    and (wand_920, a[28], b[24]) ;   // mult.v(3508)
    and (wand_951, a[29], b[23]) ;   // mult.v(3509)
    fa fa_524 (.a(wand_889), .b(wand_920), .cin(wand_951), .s(wfa_s_524), 
       .cout(wfa_cout_524));   // mult.v(3510)
    and (wand_735, a[22], b[31]) ;   // mult.v(3511)
    and (wand_766, a[23], b[30]) ;   // mult.v(3512)
    and (wand_797, a[24], b[29]) ;   // mult.v(3513)
    fa fa_525 (.a(wand_735), .b(wand_766), .cin(wand_797), .s(wfa_s_525), 
       .cout(wfa_cout_525));   // mult.v(3514)
    and (wand_828, a[25], b[28]) ;   // mult.v(3515)
    and (wand_859, a[26], b[27]) ;   // mult.v(3516)
    and (wand_890, a[27], b[26]) ;   // mult.v(3517)
    fa fa_526 (.a(wand_828), .b(wand_859), .cin(wand_890), .s(wfa_s_526), 
       .cout(wfa_cout_526));   // mult.v(3518)
    and (wand_767, a[23], b[31]) ;   // mult.v(3519)
    and (wand_798, a[24], b[30]) ;   // mult.v(3520)
    and (wand_829, a[25], b[29]) ;   // mult.v(3521)
    fa fa_527 (.a(wand_767), .b(wand_798), .cin(wand_829), .s(wfa_s_527), 
       .cout(wfa_cout_527));   // mult.v(3522)
    and (wand_6, a[0], b[6]) ;   // mult.v(3523)
    and (wand_37, a[1], b[5]) ;   // mult.v(3524)
    ha ha_24 (.a(wand_6), .b(wand_37), .s(wha_s_24), .c(wha_c_24));   // mult.v(3525)
    and (wand_7, a[0], b[7]) ;   // mult.v(3526)
    and (wand_38, a[1], b[6]) ;   // mult.v(3527)
    and (wand_69, a[2], b[5]) ;   // mult.v(3528)
    fa fa_528 (.a(wand_7), .b(wand_38), .cin(wand_69), .s(wfa_s_528), 
       .cout(wfa_cout_528));   // mult.v(3529)
    and (wand_100, a[3], b[4]) ;   // mult.v(3530)
    and (wand_131, a[4], b[3]) ;   // mult.v(3531)
    ha ha_25 (.a(wand_100), .b(wand_131), .s(wha_s_25), .c(wha_c_25));   // mult.v(3532)
    and (wand_8, a[0], b[8]) ;   // mult.v(3533)
    and (wand_39, a[1], b[7]) ;   // mult.v(3534)
    and (wand_70, a[2], b[6]) ;   // mult.v(3535)
    fa fa_529 (.a(wand_8), .b(wand_39), .cin(wand_70), .s(wfa_s_529), 
       .cout(wfa_cout_529));   // mult.v(3536)
    and (wand_101, a[3], b[5]) ;   // mult.v(3537)
    and (wand_132, a[4], b[4]) ;   // mult.v(3538)
    and (wand_163, a[5], b[3]) ;   // mult.v(3539)
    fa fa_530 (.a(wand_101), .b(wand_132), .cin(wand_163), .s(wfa_s_530), 
       .cout(wfa_cout_530));   // mult.v(3540)
    and (wand_194, a[6], b[2]) ;   // mult.v(3541)
    and (wand_225, a[7], b[1]) ;   // mult.v(3542)
    ha ha_26 (.a(wand_194), .b(wand_225), .s(wha_s_26), .c(wha_c_26));   // mult.v(3543)
    and (wand_71, a[2], b[7]) ;   // mult.v(3544)
    and (wand_102, a[3], b[6]) ;   // mult.v(3545)
    and (wand_133, a[4], b[5]) ;   // mult.v(3546)
    fa fa_531 (.a(wand_71), .b(wand_102), .cin(wand_133), .s(wfa_s_531), 
       .cout(wfa_cout_531));   // mult.v(3547)
    and (wand_164, a[5], b[4]) ;   // mult.v(3548)
    and (wand_195, a[6], b[3]) ;   // mult.v(3549)
    and (wand_226, a[7], b[2]) ;   // mult.v(3550)
    fa fa_532 (.a(wand_164), .b(wand_195), .cin(wand_226), .s(wfa_s_532), 
       .cout(wfa_cout_532));   // mult.v(3551)
    and (wand_257, a[8], b[1]) ;   // mult.v(3552)
    and (wand_288, a[9], b[0]) ;   // mult.v(3553)
    fa fa_533 (.a(wand_257), .b(wand_288), .cin(wha_s_20), .s(wfa_s_533), 
       .cout(wfa_cout_533));   // mult.v(3554)
    and (wand_165, a[5], b[5]) ;   // mult.v(3555)
    and (wand_196, a[6], b[4]) ;   // mult.v(3556)
    and (wand_227, a[7], b[3]) ;   // mult.v(3557)
    fa fa_534 (.a(wand_165), .b(wand_196), .cin(wand_227), .s(wfa_s_534), 
       .cout(wfa_cout_534));   // mult.v(3558)
    and (wand_258, a[8], b[2]) ;   // mult.v(3559)
    and (wand_289, a[9], b[1]) ;   // mult.v(3560)
    and (wand_320, a[10], b[0]) ;   // mult.v(3561)
    fa fa_535 (.a(wand_258), .b(wand_289), .cin(wand_320), .s(wfa_s_535), 
       .cout(wfa_cout_535));   // mult.v(3562)
    fa fa_536 (.a(wha_c_20), .b(wfa_s_360), .cin(wha_s_21), .s(wfa_s_536), 
       .cout(wfa_cout_536));   // mult.v(3563)
    and (wand_259, a[8], b[3]) ;   // mult.v(3564)
    and (wand_290, a[9], b[2]) ;   // mult.v(3565)
    and (wand_321, a[10], b[1]) ;   // mult.v(3566)
    fa fa_537 (.a(wand_259), .b(wand_290), .cin(wand_321), .s(wfa_s_537), 
       .cout(wfa_cout_537));   // mult.v(3567)
    and (wand_352, a[11], b[0]) ;   // mult.v(3568)
    fa fa_538 (.a(wand_352), .b(wfa_cout_360), .cin(wha_c_21), .s(wfa_s_538), 
       .cout(wfa_cout_538));   // mult.v(3569)
    fa fa_539 (.a(wfa_s_361), .b(wfa_s_362), .cin(wha_s_22), .s(wfa_s_539), 
       .cout(wfa_cout_539));   // mult.v(3570)
    and (wand_353, a[11], b[1]) ;   // mult.v(3571)
    and (wand_384, a[12], b[0]) ;   // mult.v(3572)
    fa fa_540 (.a(wand_353), .b(wand_384), .cin(wfa_cout_361), .s(wfa_s_540), 
       .cout(wfa_cout_540));   // mult.v(3573)
    fa fa_541 (.a(wfa_cout_362), .b(wha_c_22), .cin(wfa_s_363), .s(wfa_s_541), 
       .cout(wfa_cout_541));   // mult.v(3574)
    fa fa_542 (.a(wfa_s_364), .b(wfa_s_365), .cin(wha_s_23), .s(wfa_s_542), 
       .cout(wfa_cout_542));   // mult.v(3575)
    fa fa_543 (.a(wha_s_14), .b(wfa_cout_363), .cin(wfa_cout_364), .s(wfa_s_543), 
       .cout(wfa_cout_543));   // mult.v(3576)
    fa fa_544 (.a(wfa_cout_365), .b(wha_c_23), .cin(wfa_s_366), .s(wfa_s_544), 
       .cout(wfa_cout_544));   // mult.v(3577)
    fa fa_545 (.a(wfa_s_367), .b(wfa_s_368), .cin(wfa_s_369), .s(wfa_s_545), 
       .cout(wfa_cout_545));   // mult.v(3578)
    fa fa_546 (.a(wha_s_15), .b(wfa_cout_366), .cin(wfa_cout_367), .s(wfa_s_546), 
       .cout(wfa_cout_546));   // mult.v(3579)
    fa fa_547 (.a(wfa_cout_368), .b(wfa_cout_369), .cin(wfa_s_370), .s(wfa_s_547), 
       .cout(wfa_cout_547));   // mult.v(3580)
    fa fa_548 (.a(wfa_s_371), .b(wfa_s_372), .cin(wfa_s_373), .s(wfa_s_548), 
       .cout(wfa_cout_548));   // mult.v(3581)
    fa fa_549 (.a(wha_s_16), .b(wfa_cout_370), .cin(wfa_cout_371), .s(wfa_s_549), 
       .cout(wfa_cout_549));   // mult.v(3582)
    fa fa_550 (.a(wfa_cout_372), .b(wfa_cout_373), .cin(wfa_s_374), .s(wfa_s_550), 
       .cout(wfa_cout_550));   // mult.v(3583)
    fa fa_551 (.a(wfa_s_375), .b(wfa_s_376), .cin(wfa_s_377), .s(wfa_s_551), 
       .cout(wfa_cout_551));   // mult.v(3584)
    fa fa_552 (.a(wha_s_17), .b(wfa_cout_374), .cin(wfa_cout_375), .s(wfa_s_552), 
       .cout(wfa_cout_552));   // mult.v(3585)
    fa fa_553 (.a(wfa_cout_376), .b(wfa_cout_377), .cin(wfa_s_378), .s(wfa_s_553), 
       .cout(wfa_cout_553));   // mult.v(3586)
    fa fa_554 (.a(wfa_s_379), .b(wfa_s_380), .cin(wfa_s_381), .s(wfa_s_554), 
       .cout(wfa_cout_554));   // mult.v(3587)
    fa fa_555 (.a(wha_s_18), .b(wfa_cout_378), .cin(wfa_cout_379), .s(wfa_s_555), 
       .cout(wfa_cout_555));   // mult.v(3588)
    fa fa_556 (.a(wfa_cout_380), .b(wfa_cout_381), .cin(wfa_s_382), .s(wfa_s_556), 
       .cout(wfa_cout_556));   // mult.v(3589)
    fa fa_557 (.a(wfa_s_383), .b(wfa_s_384), .cin(wfa_s_385), .s(wfa_s_557), 
       .cout(wfa_cout_557));   // mult.v(3590)
    fa fa_558 (.a(wha_s_19), .b(wfa_cout_382), .cin(wfa_cout_383), .s(wfa_s_558), 
       .cout(wfa_cout_558));   // mult.v(3591)
    fa fa_559 (.a(wfa_cout_384), .b(wfa_cout_385), .cin(wfa_s_386), .s(wfa_s_559), 
       .cout(wfa_cout_559));   // mult.v(3592)
    fa fa_560 (.a(wfa_s_387), .b(wfa_s_388), .cin(wfa_s_389), .s(wfa_s_560), 
       .cout(wfa_cout_560));   // mult.v(3593)
    fa fa_561 (.a(wfa_s_188), .b(wfa_cout_386), .cin(wfa_cout_387), .s(wfa_s_561), 
       .cout(wfa_cout_561));   // mult.v(3594)
    fa fa_562 (.a(wfa_cout_388), .b(wfa_cout_389), .cin(wfa_s_390), .s(wfa_s_562), 
       .cout(wfa_cout_562));   // mult.v(3595)
    fa fa_563 (.a(wfa_s_391), .b(wfa_s_392), .cin(wfa_s_393), .s(wfa_s_563), 
       .cout(wfa_cout_563));   // mult.v(3596)
    fa fa_564 (.a(wfa_s_194), .b(wfa_cout_390), .cin(wfa_cout_391), .s(wfa_s_564), 
       .cout(wfa_cout_564));   // mult.v(3597)
    fa fa_565 (.a(wfa_cout_392), .b(wfa_cout_393), .cin(wfa_s_394), .s(wfa_s_565), 
       .cout(wfa_cout_565));   // mult.v(3598)
    fa fa_566 (.a(wfa_s_395), .b(wfa_s_396), .cin(wfa_s_397), .s(wfa_s_566), 
       .cout(wfa_cout_566));   // mult.v(3599)
    fa fa_567 (.a(wfa_s_200), .b(wfa_cout_394), .cin(wfa_cout_395), .s(wfa_s_567), 
       .cout(wfa_cout_567));   // mult.v(3600)
    fa fa_568 (.a(wfa_cout_396), .b(wfa_cout_397), .cin(wfa_s_398), .s(wfa_s_568), 
       .cout(wfa_cout_568));   // mult.v(3601)
    fa fa_569 (.a(wfa_s_399), .b(wfa_s_400), .cin(wfa_s_401), .s(wfa_s_569), 
       .cout(wfa_cout_569));   // mult.v(3602)
    fa fa_570 (.a(wfa_s_206), .b(wfa_cout_398), .cin(wfa_cout_399), .s(wfa_s_570), 
       .cout(wfa_cout_570));   // mult.v(3603)
    fa fa_571 (.a(wfa_cout_400), .b(wfa_cout_401), .cin(wfa_s_402), .s(wfa_s_571), 
       .cout(wfa_cout_571));   // mult.v(3604)
    fa fa_572 (.a(wfa_s_403), .b(wfa_s_404), .cin(wfa_s_405), .s(wfa_s_572), 
       .cout(wfa_cout_572));   // mult.v(3605)
    fa fa_573 (.a(wfa_s_212), .b(wfa_cout_402), .cin(wfa_cout_403), .s(wfa_s_573), 
       .cout(wfa_cout_573));   // mult.v(3606)
    fa fa_574 (.a(wfa_cout_404), .b(wfa_cout_405), .cin(wfa_s_406), .s(wfa_s_574), 
       .cout(wfa_cout_574));   // mult.v(3607)
    fa fa_575 (.a(wfa_s_407), .b(wfa_s_408), .cin(wfa_s_409), .s(wfa_s_575), 
       .cout(wfa_cout_575));   // mult.v(3608)
    fa fa_576 (.a(wfa_s_218), .b(wfa_cout_406), .cin(wfa_cout_407), .s(wfa_s_576), 
       .cout(wfa_cout_576));   // mult.v(3609)
    fa fa_577 (.a(wfa_cout_408), .b(wfa_cout_409), .cin(wfa_s_410), .s(wfa_s_577), 
       .cout(wfa_cout_577));   // mult.v(3610)
    fa fa_578 (.a(wfa_s_411), .b(wfa_s_412), .cin(wfa_s_413), .s(wfa_s_578), 
       .cout(wfa_cout_578));   // mult.v(3611)
    fa fa_579 (.a(wfa_s_224), .b(wfa_cout_410), .cin(wfa_cout_411), .s(wfa_s_579), 
       .cout(wfa_cout_579));   // mult.v(3612)
    fa fa_580 (.a(wfa_cout_412), .b(wfa_cout_413), .cin(wfa_s_414), .s(wfa_s_580), 
       .cout(wfa_cout_580));   // mult.v(3613)
    fa fa_581 (.a(wfa_s_415), .b(wfa_s_416), .cin(wfa_s_417), .s(wfa_s_581), 
       .cout(wfa_cout_581));   // mult.v(3614)
    fa fa_582 (.a(wfa_s_230), .b(wfa_cout_414), .cin(wfa_cout_415), .s(wfa_s_582), 
       .cout(wfa_cout_582));   // mult.v(3615)
    fa fa_583 (.a(wfa_cout_416), .b(wfa_cout_417), .cin(wfa_s_418), .s(wfa_s_583), 
       .cout(wfa_cout_583));   // mult.v(3616)
    fa fa_584 (.a(wfa_s_419), .b(wfa_s_420), .cin(wfa_s_421), .s(wfa_s_584), 
       .cout(wfa_cout_584));   // mult.v(3617)
    fa fa_585 (.a(wfa_s_236), .b(wfa_cout_418), .cin(wfa_cout_419), .s(wfa_s_585), 
       .cout(wfa_cout_585));   // mult.v(3618)
    fa fa_586 (.a(wfa_cout_420), .b(wfa_cout_421), .cin(wfa_s_422), .s(wfa_s_586), 
       .cout(wfa_cout_586));   // mult.v(3619)
    fa fa_587 (.a(wfa_s_423), .b(wfa_s_424), .cin(wfa_s_425), .s(wfa_s_587), 
       .cout(wfa_cout_587));   // mult.v(3620)
    fa fa_588 (.a(wfa_s_242), .b(wfa_cout_422), .cin(wfa_cout_423), .s(wfa_s_588), 
       .cout(wfa_cout_588));   // mult.v(3621)
    fa fa_589 (.a(wfa_cout_424), .b(wfa_cout_425), .cin(wfa_s_426), .s(wfa_s_589), 
       .cout(wfa_cout_589));   // mult.v(3622)
    fa fa_590 (.a(wfa_s_427), .b(wfa_s_428), .cin(wfa_s_429), .s(wfa_s_590), 
       .cout(wfa_cout_590));   // mult.v(3623)
    fa fa_591 (.a(wfa_s_248), .b(wfa_cout_426), .cin(wfa_cout_427), .s(wfa_s_591), 
       .cout(wfa_cout_591));   // mult.v(3624)
    fa fa_592 (.a(wfa_cout_428), .b(wfa_cout_429), .cin(wfa_s_430), .s(wfa_s_592), 
       .cout(wfa_cout_592));   // mult.v(3625)
    fa fa_593 (.a(wfa_s_431), .b(wfa_s_432), .cin(wfa_s_433), .s(wfa_s_593), 
       .cout(wfa_cout_593));   // mult.v(3626)
    fa fa_594 (.a(wfa_s_254), .b(wfa_cout_430), .cin(wfa_cout_431), .s(wfa_s_594), 
       .cout(wfa_cout_594));   // mult.v(3627)
    fa fa_595 (.a(wfa_cout_432), .b(wfa_cout_433), .cin(wfa_s_434), .s(wfa_s_595), 
       .cout(wfa_cout_595));   // mult.v(3628)
    fa fa_596 (.a(wfa_s_435), .b(wfa_s_436), .cin(wfa_s_437), .s(wfa_s_596), 
       .cout(wfa_cout_596));   // mult.v(3629)
    fa fa_597 (.a(wfa_s_260), .b(wfa_cout_434), .cin(wfa_cout_435), .s(wfa_s_597), 
       .cout(wfa_cout_597));   // mult.v(3630)
    fa fa_598 (.a(wfa_cout_436), .b(wfa_cout_437), .cin(wfa_s_438), .s(wfa_s_598), 
       .cout(wfa_cout_598));   // mult.v(3631)
    fa fa_599 (.a(wfa_s_439), .b(wfa_s_440), .cin(wfa_s_441), .s(wfa_s_599), 
       .cout(wfa_cout_599));   // mult.v(3632)
    fa fa_600 (.a(wfa_s_266), .b(wfa_cout_438), .cin(wfa_cout_439), .s(wfa_s_600), 
       .cout(wfa_cout_600));   // mult.v(3633)
    fa fa_601 (.a(wfa_cout_440), .b(wfa_cout_441), .cin(wfa_s_442), .s(wfa_s_601), 
       .cout(wfa_cout_601));   // mult.v(3634)
    fa fa_602 (.a(wfa_s_443), .b(wfa_s_444), .cin(wfa_s_445), .s(wfa_s_602), 
       .cout(wfa_cout_602));   // mult.v(3635)
    fa fa_603 (.a(wfa_s_272), .b(wfa_cout_442), .cin(wfa_cout_443), .s(wfa_s_603), 
       .cout(wfa_cout_603));   // mult.v(3636)
    fa fa_604 (.a(wfa_cout_444), .b(wfa_cout_445), .cin(wfa_s_446), .s(wfa_s_604), 
       .cout(wfa_cout_604));   // mult.v(3637)
    fa fa_605 (.a(wfa_s_447), .b(wfa_s_448), .cin(wfa_s_449), .s(wfa_s_605), 
       .cout(wfa_cout_605));   // mult.v(3638)
    fa fa_606 (.a(wfa_s_278), .b(wfa_cout_446), .cin(wfa_cout_447), .s(wfa_s_606), 
       .cout(wfa_cout_606));   // mult.v(3639)
    fa fa_607 (.a(wfa_cout_448), .b(wfa_cout_449), .cin(wfa_s_450), .s(wfa_s_607), 
       .cout(wfa_cout_607));   // mult.v(3640)
    fa fa_608 (.a(wfa_s_451), .b(wfa_s_452), .cin(wfa_s_453), .s(wfa_s_608), 
       .cout(wfa_cout_608));   // mult.v(3641)
    fa fa_609 (.a(wfa_s_284), .b(wfa_cout_450), .cin(wfa_cout_451), .s(wfa_s_609), 
       .cout(wfa_cout_609));   // mult.v(3642)
    fa fa_610 (.a(wfa_cout_452), .b(wfa_cout_453), .cin(wfa_s_454), .s(wfa_s_610), 
       .cout(wfa_cout_610));   // mult.v(3643)
    fa fa_611 (.a(wfa_s_455), .b(wfa_s_456), .cin(wfa_s_457), .s(wfa_s_611), 
       .cout(wfa_cout_611));   // mult.v(3644)
    fa fa_612 (.a(wfa_s_290), .b(wfa_cout_454), .cin(wfa_cout_455), .s(wfa_s_612), 
       .cout(wfa_cout_612));   // mult.v(3645)
    fa fa_613 (.a(wfa_cout_456), .b(wfa_cout_457), .cin(wfa_s_458), .s(wfa_s_613), 
       .cout(wfa_cout_613));   // mult.v(3646)
    fa fa_614 (.a(wfa_s_459), .b(wfa_s_460), .cin(wfa_s_461), .s(wfa_s_614), 
       .cout(wfa_cout_614));   // mult.v(3647)
    fa fa_615 (.a(wfa_s_296), .b(wfa_cout_458), .cin(wfa_cout_459), .s(wfa_s_615), 
       .cout(wfa_cout_615));   // mult.v(3648)
    fa fa_616 (.a(wfa_cout_460), .b(wfa_cout_461), .cin(wfa_s_462), .s(wfa_s_616), 
       .cout(wfa_cout_616));   // mult.v(3649)
    fa fa_617 (.a(wfa_s_463), .b(wfa_s_464), .cin(wfa_s_465), .s(wfa_s_617), 
       .cout(wfa_cout_617));   // mult.v(3650)
    fa fa_618 (.a(wfa_s_302), .b(wfa_cout_462), .cin(wfa_cout_463), .s(wfa_s_618), 
       .cout(wfa_cout_618));   // mult.v(3651)
    fa fa_619 (.a(wfa_cout_464), .b(wfa_cout_465), .cin(wfa_s_466), .s(wfa_s_619), 
       .cout(wfa_cout_619));   // mult.v(3652)
    fa fa_620 (.a(wfa_s_467), .b(wfa_s_468), .cin(wfa_s_469), .s(wfa_s_620), 
       .cout(wfa_cout_620));   // mult.v(3653)
    fa fa_621 (.a(wfa_s_308), .b(wfa_cout_466), .cin(wfa_cout_467), .s(wfa_s_621), 
       .cout(wfa_cout_621));   // mult.v(3654)
    fa fa_622 (.a(wfa_cout_468), .b(wfa_cout_469), .cin(wfa_s_470), .s(wfa_s_622), 
       .cout(wfa_cout_622));   // mult.v(3655)
    fa fa_623 (.a(wfa_s_471), .b(wfa_s_472), .cin(wfa_s_473), .s(wfa_s_623), 
       .cout(wfa_cout_623));   // mult.v(3656)
    fa fa_624 (.a(wfa_s_314), .b(wfa_cout_470), .cin(wfa_cout_471), .s(wfa_s_624), 
       .cout(wfa_cout_624));   // mult.v(3657)
    fa fa_625 (.a(wfa_cout_472), .b(wfa_cout_473), .cin(wfa_s_474), .s(wfa_s_625), 
       .cout(wfa_cout_625));   // mult.v(3658)
    fa fa_626 (.a(wfa_s_475), .b(wfa_s_476), .cin(wfa_s_477), .s(wfa_s_626), 
       .cout(wfa_cout_626));   // mult.v(3659)
    fa fa_627 (.a(wfa_s_320), .b(wfa_cout_474), .cin(wfa_cout_475), .s(wfa_s_627), 
       .cout(wfa_cout_627));   // mult.v(3660)
    fa fa_628 (.a(wfa_cout_476), .b(wfa_cout_477), .cin(wfa_s_478), .s(wfa_s_628), 
       .cout(wfa_cout_628));   // mult.v(3661)
    fa fa_629 (.a(wfa_s_479), .b(wfa_s_480), .cin(wfa_s_481), .s(wfa_s_629), 
       .cout(wfa_cout_629));   // mult.v(3662)
    fa fa_630 (.a(wfa_s_326), .b(wfa_cout_478), .cin(wfa_cout_479), .s(wfa_s_630), 
       .cout(wfa_cout_630));   // mult.v(3663)
    fa fa_631 (.a(wfa_cout_480), .b(wfa_cout_481), .cin(wfa_s_482), .s(wfa_s_631), 
       .cout(wfa_cout_631));   // mult.v(3664)
    fa fa_632 (.a(wfa_s_483), .b(wfa_s_484), .cin(wfa_s_485), .s(wfa_s_632), 
       .cout(wfa_cout_632));   // mult.v(3665)
    fa fa_633 (.a(wfa_s_332), .b(wfa_cout_482), .cin(wfa_cout_483), .s(wfa_s_633), 
       .cout(wfa_cout_633));   // mult.v(3666)
    fa fa_634 (.a(wfa_cout_484), .b(wfa_cout_485), .cin(wfa_s_486), .s(wfa_s_634), 
       .cout(wfa_cout_634));   // mult.v(3667)
    fa fa_635 (.a(wfa_s_487), .b(wfa_s_488), .cin(wfa_s_489), .s(wfa_s_635), 
       .cout(wfa_cout_635));   // mult.v(3668)
    fa fa_636 (.a(wfa_s_338), .b(wfa_cout_486), .cin(wfa_cout_487), .s(wfa_s_636), 
       .cout(wfa_cout_636));   // mult.v(3669)
    fa fa_637 (.a(wfa_cout_488), .b(wfa_cout_489), .cin(wfa_s_490), .s(wfa_s_637), 
       .cout(wfa_cout_637));   // mult.v(3670)
    fa fa_638 (.a(wfa_s_491), .b(wfa_s_492), .cin(wfa_s_493), .s(wfa_s_638), 
       .cout(wfa_cout_638));   // mult.v(3671)
    fa fa_639 (.a(wfa_s_344), .b(wfa_cout_490), .cin(wfa_cout_491), .s(wfa_s_639), 
       .cout(wfa_cout_639));   // mult.v(3672)
    fa fa_640 (.a(wfa_cout_492), .b(wfa_cout_493), .cin(wfa_s_494), .s(wfa_s_640), 
       .cout(wfa_cout_640));   // mult.v(3673)
    fa fa_641 (.a(wfa_s_495), .b(wfa_s_496), .cin(wfa_s_497), .s(wfa_s_641), 
       .cout(wfa_cout_641));   // mult.v(3674)
    fa fa_642 (.a(wfa_s_349), .b(wfa_cout_494), .cin(wfa_cout_495), .s(wfa_s_642), 
       .cout(wfa_cout_642));   // mult.v(3675)
    fa fa_643 (.a(wfa_cout_496), .b(wfa_cout_497), .cin(wfa_s_498), .s(wfa_s_643), 
       .cout(wfa_cout_643));   // mult.v(3676)
    fa fa_644 (.a(wfa_s_499), .b(wfa_s_500), .cin(wfa_s_501), .s(wfa_s_644), 
       .cout(wfa_cout_644));   // mult.v(3677)
    fa fa_645 (.a(wfa_s_353), .b(wfa_cout_498), .cin(wfa_cout_499), .s(wfa_s_645), 
       .cout(wfa_cout_645));   // mult.v(3678)
    fa fa_646 (.a(wfa_cout_500), .b(wfa_cout_501), .cin(wfa_s_502), .s(wfa_s_646), 
       .cout(wfa_cout_646));   // mult.v(3679)
    fa fa_647 (.a(wfa_s_503), .b(wfa_s_504), .cin(wfa_s_505), .s(wfa_s_647), 
       .cout(wfa_cout_647));   // mult.v(3680)
    fa fa_648 (.a(wfa_s_356), .b(wfa_cout_502), .cin(wfa_cout_503), .s(wfa_s_648), 
       .cout(wfa_cout_648));   // mult.v(3681)
    fa fa_649 (.a(wfa_cout_504), .b(wfa_cout_505), .cin(wfa_s_506), .s(wfa_s_649), 
       .cout(wfa_cout_649));   // mult.v(3682)
    fa fa_650 (.a(wfa_s_507), .b(wfa_s_508), .cin(wfa_s_509), .s(wfa_s_650), 
       .cout(wfa_cout_650));   // mult.v(3683)
    fa fa_651 (.a(wfa_s_358), .b(wfa_cout_506), .cin(wfa_cout_507), .s(wfa_s_651), 
       .cout(wfa_cout_651));   // mult.v(3684)
    fa fa_652 (.a(wfa_cout_508), .b(wfa_cout_509), .cin(wfa_s_510), .s(wfa_s_652), 
       .cout(wfa_cout_652));   // mult.v(3685)
    fa fa_653 (.a(wfa_s_511), .b(wfa_s_512), .cin(wfa_s_513), .s(wfa_s_653), 
       .cout(wfa_cout_653));   // mult.v(3686)
    fa fa_654 (.a(wfa_s_359), .b(wfa_cout_510), .cin(wfa_cout_511), .s(wfa_s_654), 
       .cout(wfa_cout_654));   // mult.v(3687)
    fa fa_655 (.a(wfa_cout_512), .b(wfa_cout_513), .cin(wfa_s_514), .s(wfa_s_655), 
       .cout(wfa_cout_655));   // mult.v(3688)
    fa fa_656 (.a(wfa_s_515), .b(wfa_s_516), .cin(wfa_s_517), .s(wfa_s_656), 
       .cout(wfa_cout_656));   // mult.v(3689)
    fa fa_657 (.a(wfa_cout_359), .b(wfa_cout_514), .cin(wfa_cout_515), 
       .s(wfa_s_657), .cout(wfa_cout_657));   // mult.v(3690)
    fa fa_658 (.a(wfa_cout_516), .b(wfa_cout_517), .cin(wfa_s_518), .s(wfa_s_658), 
       .cout(wfa_cout_658));   // mult.v(3691)
    fa fa_659 (.a(wfa_s_519), .b(wfa_s_520), .cin(wfa_s_521), .s(wfa_s_659), 
       .cout(wfa_cout_659));   // mult.v(3692)
    and (wand_982, a[30], b[22]) ;   // mult.v(3693)
    and (wand_1013, a[31], b[21]) ;   // mult.v(3694)
    fa fa_660 (.a(wand_982), .b(wand_1013), .cin(wfa_cout_518), .s(wfa_s_660), 
       .cout(wfa_cout_660));   // mult.v(3695)
    fa fa_661 (.a(wfa_cout_519), .b(wfa_cout_520), .cin(wfa_cout_521), 
       .s(wfa_s_661), .cout(wfa_cout_661));   // mult.v(3696)
    fa fa_662 (.a(wfa_s_522), .b(wfa_s_523), .cin(wfa_s_524), .s(wfa_s_662), 
       .cout(wfa_cout_662));   // mult.v(3697)
    and (wand_921, a[28], b[25]) ;   // mult.v(3698)
    and (wand_952, a[29], b[24]) ;   // mult.v(3699)
    and (wand_983, a[30], b[23]) ;   // mult.v(3700)
    fa fa_663 (.a(wand_921), .b(wand_952), .cin(wand_983), .s(wfa_s_663), 
       .cout(wfa_cout_663));   // mult.v(3701)
    and (wand_1014, a[31], b[22]) ;   // mult.v(3702)
    fa fa_664 (.a(wand_1014), .b(wfa_cout_522), .cin(wfa_cout_523), .s(wfa_s_664), 
       .cout(wfa_cout_664));   // mult.v(3703)
    fa fa_665 (.a(wfa_cout_524), .b(wfa_s_525), .cin(wfa_s_526), .s(wfa_s_665), 
       .cout(wfa_cout_665));   // mult.v(3704)
    and (wand_860, a[26], b[28]) ;   // mult.v(3705)
    and (wand_891, a[27], b[27]) ;   // mult.v(3706)
    and (wand_922, a[28], b[26]) ;   // mult.v(3707)
    fa fa_666 (.a(wand_860), .b(wand_891), .cin(wand_922), .s(wfa_s_666), 
       .cout(wfa_cout_666));   // mult.v(3708)
    and (wand_953, a[29], b[25]) ;   // mult.v(3709)
    and (wand_984, a[30], b[24]) ;   // mult.v(3710)
    and (wand_1015, a[31], b[23]) ;   // mult.v(3711)
    fa fa_667 (.a(wand_953), .b(wand_984), .cin(wand_1015), .s(wfa_s_667), 
       .cout(wfa_cout_667));   // mult.v(3712)
    fa fa_668 (.a(wfa_cout_525), .b(wfa_cout_526), .cin(wfa_s_527), .s(wfa_s_668), 
       .cout(wfa_cout_668));   // mult.v(3713)
    and (wand_799, a[24], b[31]) ;   // mult.v(3714)
    and (wand_830, a[25], b[30]) ;   // mult.v(3715)
    and (wand_861, a[26], b[29]) ;   // mult.v(3716)
    fa fa_669 (.a(wand_799), .b(wand_830), .cin(wand_861), .s(wfa_s_669), 
       .cout(wfa_cout_669));   // mult.v(3717)
    and (wand_892, a[27], b[28]) ;   // mult.v(3718)
    and (wand_923, a[28], b[27]) ;   // mult.v(3719)
    and (wand_954, a[29], b[26]) ;   // mult.v(3720)
    fa fa_670 (.a(wand_892), .b(wand_923), .cin(wand_954), .s(wfa_s_670), 
       .cout(wfa_cout_670));   // mult.v(3721)
    and (wand_985, a[30], b[25]) ;   // mult.v(3722)
    and (wand_1016, a[31], b[24]) ;   // mult.v(3723)
    fa fa_671 (.a(wand_985), .b(wand_1016), .cin(wfa_cout_527), .s(wfa_s_671), 
       .cout(wfa_cout_671));   // mult.v(3724)
    and (wand_831, a[25], b[31]) ;   // mult.v(3725)
    and (wand_862, a[26], b[30]) ;   // mult.v(3726)
    and (wand_893, a[27], b[29]) ;   // mult.v(3727)
    fa fa_672 (.a(wand_831), .b(wand_862), .cin(wand_893), .s(wfa_s_672), 
       .cout(wfa_cout_672));   // mult.v(3728)
    and (wand_924, a[28], b[28]) ;   // mult.v(3729)
    and (wand_955, a[29], b[27]) ;   // mult.v(3730)
    and (wand_986, a[30], b[26]) ;   // mult.v(3731)
    fa fa_673 (.a(wand_924), .b(wand_955), .cin(wand_986), .s(wfa_s_673), 
       .cout(wfa_cout_673));   // mult.v(3732)
    and (wand_863, a[26], b[31]) ;   // mult.v(3733)
    and (wand_894, a[27], b[30]) ;   // mult.v(3734)
    and (wand_925, a[28], b[29]) ;   // mult.v(3735)
    fa fa_674 (.a(wand_863), .b(wand_894), .cin(wand_925), .s(wfa_s_674), 
       .cout(wfa_cout_674));   // mult.v(3736)
    and (wand_4, a[0], b[4]) ;   // mult.v(3737)
    and (wand_35, a[1], b[3]) ;   // mult.v(3738)
    ha ha_27 (.a(wand_4), .b(wand_35), .s(wha_s_27), .c(wha_c_27));   // mult.v(3739)
    and (wand_5, a[0], b[5]) ;   // mult.v(3740)
    and (wand_36, a[1], b[4]) ;   // mult.v(3741)
    and (wand_67, a[2], b[3]) ;   // mult.v(3742)
    fa fa_675 (.a(wand_5), .b(wand_36), .cin(wand_67), .s(wfa_s_675), 
       .cout(wfa_cout_675));   // mult.v(3743)
    and (wand_98, a[3], b[2]) ;   // mult.v(3744)
    and (wand_129, a[4], b[1]) ;   // mult.v(3745)
    ha ha_28 (.a(wand_98), .b(wand_129), .s(wha_s_28), .c(wha_c_28));   // mult.v(3746)
    and (wand_68, a[2], b[4]) ;   // mult.v(3747)
    and (wand_99, a[3], b[3]) ;   // mult.v(3748)
    and (wand_130, a[4], b[2]) ;   // mult.v(3749)
    fa fa_676 (.a(wand_68), .b(wand_99), .cin(wand_130), .s(wfa_s_676), 
       .cout(wfa_cout_676));   // mult.v(3750)
    and (wand_161, a[5], b[1]) ;   // mult.v(3751)
    and (wand_192, a[6], b[0]) ;   // mult.v(3752)
    fa fa_677 (.a(wand_161), .b(wand_192), .cin(wha_s_24), .s(wfa_s_677), 
       .cout(wfa_cout_677));   // mult.v(3753)
    and (wand_162, a[5], b[2]) ;   // mult.v(3754)
    and (wand_193, a[6], b[1]) ;   // mult.v(3755)
    and (wand_224, a[7], b[0]) ;   // mult.v(3756)
    fa fa_678 (.a(wand_162), .b(wand_193), .cin(wand_224), .s(wfa_s_678), 
       .cout(wfa_cout_678));   // mult.v(3757)
    fa fa_679 (.a(wha_c_24), .b(wfa_s_528), .cin(wha_s_25), .s(wfa_s_679), 
       .cout(wfa_cout_679));   // mult.v(3758)
    and (wand_256, a[8], b[0]) ;   // mult.v(3759)
    fa fa_680 (.a(wand_256), .b(wfa_cout_528), .cin(wha_c_25), .s(wfa_s_680), 
       .cout(wfa_cout_680));   // mult.v(3760)
    fa fa_681 (.a(wfa_s_529), .b(wfa_s_530), .cin(wha_s_26), .s(wfa_s_681), 
       .cout(wfa_cout_681));   // mult.v(3761)
    fa fa_682 (.a(wfa_cout_529), .b(wfa_cout_530), .cin(wha_c_26), .s(wfa_s_682), 
       .cout(wfa_cout_682));   // mult.v(3762)
    fa fa_683 (.a(wfa_s_531), .b(wfa_s_532), .cin(wfa_s_533), .s(wfa_s_683), 
       .cout(wfa_cout_683));   // mult.v(3763)
    fa fa_684 (.a(wfa_cout_531), .b(wfa_cout_532), .cin(wfa_cout_533), 
       .s(wfa_s_684), .cout(wfa_cout_684));   // mult.v(3764)
    fa fa_685 (.a(wfa_s_534), .b(wfa_s_535), .cin(wfa_s_536), .s(wfa_s_685), 
       .cout(wfa_cout_685));   // mult.v(3765)
    fa fa_686 (.a(wfa_cout_534), .b(wfa_cout_535), .cin(wfa_cout_536), 
       .s(wfa_s_686), .cout(wfa_cout_686));   // mult.v(3766)
    fa fa_687 (.a(wfa_s_537), .b(wfa_s_538), .cin(wfa_s_539), .s(wfa_s_687), 
       .cout(wfa_cout_687));   // mult.v(3767)
    fa fa_688 (.a(wfa_cout_537), .b(wfa_cout_538), .cin(wfa_cout_539), 
       .s(wfa_s_688), .cout(wfa_cout_688));   // mult.v(3768)
    fa fa_689 (.a(wfa_s_540), .b(wfa_s_541), .cin(wfa_s_542), .s(wfa_s_689), 
       .cout(wfa_cout_689));   // mult.v(3769)
    fa fa_690 (.a(wfa_cout_540), .b(wfa_cout_541), .cin(wfa_cout_542), 
       .s(wfa_s_690), .cout(wfa_cout_690));   // mult.v(3770)
    fa fa_691 (.a(wfa_s_543), .b(wfa_s_544), .cin(wfa_s_545), .s(wfa_s_691), 
       .cout(wfa_cout_691));   // mult.v(3771)
    fa fa_692 (.a(wfa_cout_543), .b(wfa_cout_544), .cin(wfa_cout_545), 
       .s(wfa_s_692), .cout(wfa_cout_692));   // mult.v(3772)
    fa fa_693 (.a(wfa_s_546), .b(wfa_s_547), .cin(wfa_s_548), .s(wfa_s_693), 
       .cout(wfa_cout_693));   // mult.v(3773)
    fa fa_694 (.a(wfa_cout_546), .b(wfa_cout_547), .cin(wfa_cout_548), 
       .s(wfa_s_694), .cout(wfa_cout_694));   // mult.v(3774)
    fa fa_695 (.a(wfa_s_549), .b(wfa_s_550), .cin(wfa_s_551), .s(wfa_s_695), 
       .cout(wfa_cout_695));   // mult.v(3775)
    fa fa_696 (.a(wfa_cout_549), .b(wfa_cout_550), .cin(wfa_cout_551), 
       .s(wfa_s_696), .cout(wfa_cout_696));   // mult.v(3776)
    fa fa_697 (.a(wfa_s_552), .b(wfa_s_553), .cin(wfa_s_554), .s(wfa_s_697), 
       .cout(wfa_cout_697));   // mult.v(3777)
    fa fa_698 (.a(wfa_cout_552), .b(wfa_cout_553), .cin(wfa_cout_554), 
       .s(wfa_s_698), .cout(wfa_cout_698));   // mult.v(3778)
    fa fa_699 (.a(wfa_s_555), .b(wfa_s_556), .cin(wfa_s_557), .s(wfa_s_699), 
       .cout(wfa_cout_699));   // mult.v(3779)
    fa fa_700 (.a(wfa_cout_555), .b(wfa_cout_556), .cin(wfa_cout_557), 
       .s(wfa_s_700), .cout(wfa_cout_700));   // mult.v(3780)
    fa fa_701 (.a(wfa_s_558), .b(wfa_s_559), .cin(wfa_s_560), .s(wfa_s_701), 
       .cout(wfa_cout_701));   // mult.v(3781)
    fa fa_702 (.a(wfa_cout_558), .b(wfa_cout_559), .cin(wfa_cout_560), 
       .s(wfa_s_702), .cout(wfa_cout_702));   // mult.v(3782)
    fa fa_703 (.a(wfa_s_561), .b(wfa_s_562), .cin(wfa_s_563), .s(wfa_s_703), 
       .cout(wfa_cout_703));   // mult.v(3783)
    fa fa_704 (.a(wfa_cout_561), .b(wfa_cout_562), .cin(wfa_cout_563), 
       .s(wfa_s_704), .cout(wfa_cout_704));   // mult.v(3784)
    fa fa_705 (.a(wfa_s_564), .b(wfa_s_565), .cin(wfa_s_566), .s(wfa_s_705), 
       .cout(wfa_cout_705));   // mult.v(3785)
    fa fa_706 (.a(wfa_cout_564), .b(wfa_cout_565), .cin(wfa_cout_566), 
       .s(wfa_s_706), .cout(wfa_cout_706));   // mult.v(3786)
    fa fa_707 (.a(wfa_s_567), .b(wfa_s_568), .cin(wfa_s_569), .s(wfa_s_707), 
       .cout(wfa_cout_707));   // mult.v(3787)
    fa fa_708 (.a(wfa_cout_567), .b(wfa_cout_568), .cin(wfa_cout_569), 
       .s(wfa_s_708), .cout(wfa_cout_708));   // mult.v(3788)
    fa fa_709 (.a(wfa_s_570), .b(wfa_s_571), .cin(wfa_s_572), .s(wfa_s_709), 
       .cout(wfa_cout_709));   // mult.v(3789)
    fa fa_710 (.a(wfa_cout_570), .b(wfa_cout_571), .cin(wfa_cout_572), 
       .s(wfa_s_710), .cout(wfa_cout_710));   // mult.v(3790)
    fa fa_711 (.a(wfa_s_573), .b(wfa_s_574), .cin(wfa_s_575), .s(wfa_s_711), 
       .cout(wfa_cout_711));   // mult.v(3791)
    fa fa_712 (.a(wfa_cout_573), .b(wfa_cout_574), .cin(wfa_cout_575), 
       .s(wfa_s_712), .cout(wfa_cout_712));   // mult.v(3792)
    fa fa_713 (.a(wfa_s_576), .b(wfa_s_577), .cin(wfa_s_578), .s(wfa_s_713), 
       .cout(wfa_cout_713));   // mult.v(3793)
    fa fa_714 (.a(wfa_cout_576), .b(wfa_cout_577), .cin(wfa_cout_578), 
       .s(wfa_s_714), .cout(wfa_cout_714));   // mult.v(3794)
    fa fa_715 (.a(wfa_s_579), .b(wfa_s_580), .cin(wfa_s_581), .s(wfa_s_715), 
       .cout(wfa_cout_715));   // mult.v(3795)
    fa fa_716 (.a(wfa_cout_579), .b(wfa_cout_580), .cin(wfa_cout_581), 
       .s(wfa_s_716), .cout(wfa_cout_716));   // mult.v(3796)
    fa fa_717 (.a(wfa_s_582), .b(wfa_s_583), .cin(wfa_s_584), .s(wfa_s_717), 
       .cout(wfa_cout_717));   // mult.v(3797)
    fa fa_718 (.a(wfa_cout_582), .b(wfa_cout_583), .cin(wfa_cout_584), 
       .s(wfa_s_718), .cout(wfa_cout_718));   // mult.v(3798)
    fa fa_719 (.a(wfa_s_585), .b(wfa_s_586), .cin(wfa_s_587), .s(wfa_s_719), 
       .cout(wfa_cout_719));   // mult.v(3799)
    fa fa_720 (.a(wfa_cout_585), .b(wfa_cout_586), .cin(wfa_cout_587), 
       .s(wfa_s_720), .cout(wfa_cout_720));   // mult.v(3800)
    fa fa_721 (.a(wfa_s_588), .b(wfa_s_589), .cin(wfa_s_590), .s(wfa_s_721), 
       .cout(wfa_cout_721));   // mult.v(3801)
    fa fa_722 (.a(wfa_cout_588), .b(wfa_cout_589), .cin(wfa_cout_590), 
       .s(wfa_s_722), .cout(wfa_cout_722));   // mult.v(3802)
    fa fa_723 (.a(wfa_s_591), .b(wfa_s_592), .cin(wfa_s_593), .s(wfa_s_723), 
       .cout(wfa_cout_723));   // mult.v(3803)
    fa fa_724 (.a(wfa_cout_591), .b(wfa_cout_592), .cin(wfa_cout_593), 
       .s(wfa_s_724), .cout(wfa_cout_724));   // mult.v(3804)
    fa fa_725 (.a(wfa_s_594), .b(wfa_s_595), .cin(wfa_s_596), .s(wfa_s_725), 
       .cout(wfa_cout_725));   // mult.v(3805)
    fa fa_726 (.a(wfa_cout_594), .b(wfa_cout_595), .cin(wfa_cout_596), 
       .s(wfa_s_726), .cout(wfa_cout_726));   // mult.v(3806)
    fa fa_727 (.a(wfa_s_597), .b(wfa_s_598), .cin(wfa_s_599), .s(wfa_s_727), 
       .cout(wfa_cout_727));   // mult.v(3807)
    fa fa_728 (.a(wfa_cout_597), .b(wfa_cout_598), .cin(wfa_cout_599), 
       .s(wfa_s_728), .cout(wfa_cout_728));   // mult.v(3808)
    fa fa_729 (.a(wfa_s_600), .b(wfa_s_601), .cin(wfa_s_602), .s(wfa_s_729), 
       .cout(wfa_cout_729));   // mult.v(3809)
    fa fa_730 (.a(wfa_cout_600), .b(wfa_cout_601), .cin(wfa_cout_602), 
       .s(wfa_s_730), .cout(wfa_cout_730));   // mult.v(3810)
    fa fa_731 (.a(wfa_s_603), .b(wfa_s_604), .cin(wfa_s_605), .s(wfa_s_731), 
       .cout(wfa_cout_731));   // mult.v(3811)
    fa fa_732 (.a(wfa_cout_603), .b(wfa_cout_604), .cin(wfa_cout_605), 
       .s(wfa_s_732), .cout(wfa_cout_732));   // mult.v(3812)
    fa fa_733 (.a(wfa_s_606), .b(wfa_s_607), .cin(wfa_s_608), .s(wfa_s_733), 
       .cout(wfa_cout_733));   // mult.v(3813)
    fa fa_734 (.a(wfa_cout_606), .b(wfa_cout_607), .cin(wfa_cout_608), 
       .s(wfa_s_734), .cout(wfa_cout_734));   // mult.v(3814)
    fa fa_735 (.a(wfa_s_609), .b(wfa_s_610), .cin(wfa_s_611), .s(wfa_s_735), 
       .cout(wfa_cout_735));   // mult.v(3815)
    fa fa_736 (.a(wfa_cout_609), .b(wfa_cout_610), .cin(wfa_cout_611), 
       .s(wfa_s_736), .cout(wfa_cout_736));   // mult.v(3816)
    fa fa_737 (.a(wfa_s_612), .b(wfa_s_613), .cin(wfa_s_614), .s(wfa_s_737), 
       .cout(wfa_cout_737));   // mult.v(3817)
    fa fa_738 (.a(wfa_cout_612), .b(wfa_cout_613), .cin(wfa_cout_614), 
       .s(wfa_s_738), .cout(wfa_cout_738));   // mult.v(3818)
    fa fa_739 (.a(wfa_s_615), .b(wfa_s_616), .cin(wfa_s_617), .s(wfa_s_739), 
       .cout(wfa_cout_739));   // mult.v(3819)
    fa fa_740 (.a(wfa_cout_615), .b(wfa_cout_616), .cin(wfa_cout_617), 
       .s(wfa_s_740), .cout(wfa_cout_740));   // mult.v(3820)
    fa fa_741 (.a(wfa_s_618), .b(wfa_s_619), .cin(wfa_s_620), .s(wfa_s_741), 
       .cout(wfa_cout_741));   // mult.v(3821)
    fa fa_742 (.a(wfa_cout_618), .b(wfa_cout_619), .cin(wfa_cout_620), 
       .s(wfa_s_742), .cout(wfa_cout_742));   // mult.v(3822)
    fa fa_743 (.a(wfa_s_621), .b(wfa_s_622), .cin(wfa_s_623), .s(wfa_s_743), 
       .cout(wfa_cout_743));   // mult.v(3823)
    fa fa_744 (.a(wfa_cout_621), .b(wfa_cout_622), .cin(wfa_cout_623), 
       .s(wfa_s_744), .cout(wfa_cout_744));   // mult.v(3824)
    fa fa_745 (.a(wfa_s_624), .b(wfa_s_625), .cin(wfa_s_626), .s(wfa_s_745), 
       .cout(wfa_cout_745));   // mult.v(3825)
    fa fa_746 (.a(wfa_cout_624), .b(wfa_cout_625), .cin(wfa_cout_626), 
       .s(wfa_s_746), .cout(wfa_cout_746));   // mult.v(3826)
    fa fa_747 (.a(wfa_s_627), .b(wfa_s_628), .cin(wfa_s_629), .s(wfa_s_747), 
       .cout(wfa_cout_747));   // mult.v(3827)
    fa fa_748 (.a(wfa_cout_627), .b(wfa_cout_628), .cin(wfa_cout_629), 
       .s(wfa_s_748), .cout(wfa_cout_748));   // mult.v(3828)
    fa fa_749 (.a(wfa_s_630), .b(wfa_s_631), .cin(wfa_s_632), .s(wfa_s_749), 
       .cout(wfa_cout_749));   // mult.v(3829)
    fa fa_750 (.a(wfa_cout_630), .b(wfa_cout_631), .cin(wfa_cout_632), 
       .s(wfa_s_750), .cout(wfa_cout_750));   // mult.v(3830)
    fa fa_751 (.a(wfa_s_633), .b(wfa_s_634), .cin(wfa_s_635), .s(wfa_s_751), 
       .cout(wfa_cout_751));   // mult.v(3831)
    fa fa_752 (.a(wfa_cout_633), .b(wfa_cout_634), .cin(wfa_cout_635), 
       .s(wfa_s_752), .cout(wfa_cout_752));   // mult.v(3832)
    fa fa_753 (.a(wfa_s_636), .b(wfa_s_637), .cin(wfa_s_638), .s(wfa_s_753), 
       .cout(wfa_cout_753));   // mult.v(3833)
    fa fa_754 (.a(wfa_cout_636), .b(wfa_cout_637), .cin(wfa_cout_638), 
       .s(wfa_s_754), .cout(wfa_cout_754));   // mult.v(3834)
    fa fa_755 (.a(wfa_s_639), .b(wfa_s_640), .cin(wfa_s_641), .s(wfa_s_755), 
       .cout(wfa_cout_755));   // mult.v(3835)
    fa fa_756 (.a(wfa_cout_639), .b(wfa_cout_640), .cin(wfa_cout_641), 
       .s(wfa_s_756), .cout(wfa_cout_756));   // mult.v(3836)
    fa fa_757 (.a(wfa_s_642), .b(wfa_s_643), .cin(wfa_s_644), .s(wfa_s_757), 
       .cout(wfa_cout_757));   // mult.v(3837)
    fa fa_758 (.a(wfa_cout_642), .b(wfa_cout_643), .cin(wfa_cout_644), 
       .s(wfa_s_758), .cout(wfa_cout_758));   // mult.v(3838)
    fa fa_759 (.a(wfa_s_645), .b(wfa_s_646), .cin(wfa_s_647), .s(wfa_s_759), 
       .cout(wfa_cout_759));   // mult.v(3839)
    fa fa_760 (.a(wfa_cout_645), .b(wfa_cout_646), .cin(wfa_cout_647), 
       .s(wfa_s_760), .cout(wfa_cout_760));   // mult.v(3840)
    fa fa_761 (.a(wfa_s_648), .b(wfa_s_649), .cin(wfa_s_650), .s(wfa_s_761), 
       .cout(wfa_cout_761));   // mult.v(3841)
    fa fa_762 (.a(wfa_cout_648), .b(wfa_cout_649), .cin(wfa_cout_650), 
       .s(wfa_s_762), .cout(wfa_cout_762));   // mult.v(3842)
    fa fa_763 (.a(wfa_s_651), .b(wfa_s_652), .cin(wfa_s_653), .s(wfa_s_763), 
       .cout(wfa_cout_763));   // mult.v(3843)
    fa fa_764 (.a(wfa_cout_651), .b(wfa_cout_652), .cin(wfa_cout_653), 
       .s(wfa_s_764), .cout(wfa_cout_764));   // mult.v(3844)
    fa fa_765 (.a(wfa_s_654), .b(wfa_s_655), .cin(wfa_s_656), .s(wfa_s_765), 
       .cout(wfa_cout_765));   // mult.v(3845)
    fa fa_766 (.a(wfa_cout_654), .b(wfa_cout_655), .cin(wfa_cout_656), 
       .s(wfa_s_766), .cout(wfa_cout_766));   // mult.v(3846)
    fa fa_767 (.a(wfa_s_657), .b(wfa_s_658), .cin(wfa_s_659), .s(wfa_s_767), 
       .cout(wfa_cout_767));   // mult.v(3847)
    fa fa_768 (.a(wfa_cout_657), .b(wfa_cout_658), .cin(wfa_cout_659), 
       .s(wfa_s_768), .cout(wfa_cout_768));   // mult.v(3848)
    fa fa_769 (.a(wfa_s_660), .b(wfa_s_661), .cin(wfa_s_662), .s(wfa_s_769), 
       .cout(wfa_cout_769));   // mult.v(3849)
    fa fa_770 (.a(wfa_cout_660), .b(wfa_cout_661), .cin(wfa_cout_662), 
       .s(wfa_s_770), .cout(wfa_cout_770));   // mult.v(3850)
    fa fa_771 (.a(wfa_s_663), .b(wfa_s_664), .cin(wfa_s_665), .s(wfa_s_771), 
       .cout(wfa_cout_771));   // mult.v(3851)
    fa fa_772 (.a(wfa_cout_663), .b(wfa_cout_664), .cin(wfa_cout_665), 
       .s(wfa_s_772), .cout(wfa_cout_772));   // mult.v(3852)
    fa fa_773 (.a(wfa_s_666), .b(wfa_s_667), .cin(wfa_s_668), .s(wfa_s_773), 
       .cout(wfa_cout_773));   // mult.v(3853)
    fa fa_774 (.a(wfa_cout_666), .b(wfa_cout_667), .cin(wfa_cout_668), 
       .s(wfa_s_774), .cout(wfa_cout_774));   // mult.v(3854)
    fa fa_775 (.a(wfa_s_669), .b(wfa_s_670), .cin(wfa_s_671), .s(wfa_s_775), 
       .cout(wfa_cout_775));   // mult.v(3855)
    and (wand_1017, a[31], b[25]) ;   // mult.v(3856)
    fa fa_776 (.a(wand_1017), .b(wfa_cout_669), .cin(wfa_cout_670), .s(wfa_s_776), 
       .cout(wfa_cout_776));   // mult.v(3857)
    fa fa_777 (.a(wfa_cout_671), .b(wfa_s_672), .cin(wfa_s_673), .s(wfa_s_777), 
       .cout(wfa_cout_777));   // mult.v(3858)
    and (wand_956, a[29], b[28]) ;   // mult.v(3859)
    and (wand_987, a[30], b[27]) ;   // mult.v(3860)
    and (wand_1018, a[31], b[26]) ;   // mult.v(3861)
    fa fa_778 (.a(wand_956), .b(wand_987), .cin(wand_1018), .s(wfa_s_778), 
       .cout(wfa_cout_778));   // mult.v(3862)
    fa fa_779 (.a(wfa_cout_672), .b(wfa_cout_673), .cin(wfa_s_674), .s(wfa_s_779), 
       .cout(wfa_cout_779));   // mult.v(3863)
    and (wand_895, a[27], b[31]) ;   // mult.v(3864)
    and (wand_926, a[28], b[30]) ;   // mult.v(3865)
    and (wand_957, a[29], b[29]) ;   // mult.v(3866)
    fa fa_780 (.a(wand_895), .b(wand_926), .cin(wand_957), .s(wfa_s_780), 
       .cout(wfa_cout_780));   // mult.v(3867)
    and (wand_988, a[30], b[28]) ;   // mult.v(3868)
    and (wand_1019, a[31], b[27]) ;   // mult.v(3869)
    fa fa_781 (.a(wand_988), .b(wand_1019), .cin(wfa_cout_674), .s(wfa_s_781), 
       .cout(wfa_cout_781));   // mult.v(3870)
    and (wand_927, a[28], b[31]) ;   // mult.v(3871)
    and (wand_958, a[29], b[30]) ;   // mult.v(3872)
    and (wand_989, a[30], b[29]) ;   // mult.v(3873)
    fa fa_782 (.a(wand_927), .b(wand_958), .cin(wand_989), .s(wfa_s_782), 
       .cout(wfa_cout_782));   // mult.v(3874)
    and (wand_3, a[0], b[3]) ;   // mult.v(3875)
    and (wand_34, a[1], b[2]) ;   // mult.v(3876)
    ha ha_29 (.a(wand_3), .b(wand_34), .s(wha_s_29), .c(wha_c_29));   // mult.v(3877)
    and (wand_66, a[2], b[2]) ;   // mult.v(3878)
    and (wand_97, a[3], b[1]) ;   // mult.v(3879)
    and (wand_128, a[4], b[0]) ;   // mult.v(3880)
    fa fa_783 (.a(wand_66), .b(wand_97), .cin(wand_128), .s(wfa_s_783), 
       .cout(wfa_cout_783));   // mult.v(3881)
    and (wand_160, a[5], b[0]) ;   // mult.v(3882)
    fa fa_784 (.a(wand_160), .b(wha_c_27), .cin(wfa_s_675), .s(wfa_s_784), 
       .cout(wfa_cout_784));   // mult.v(3883)
    fa fa_785 (.a(wfa_cout_675), .b(wha_c_28), .cin(wfa_s_676), .s(wfa_s_785), 
       .cout(wfa_cout_785));   // mult.v(3884)
    fa fa_786 (.a(wfa_cout_676), .b(wfa_cout_677), .cin(wfa_s_678), .s(wfa_s_786), 
       .cout(wfa_cout_786));   // mult.v(3885)
    fa fa_787 (.a(wfa_cout_678), .b(wfa_cout_679), .cin(wfa_s_680), .s(wfa_s_787), 
       .cout(wfa_cout_787));   // mult.v(3886)
    fa fa_788 (.a(wfa_cout_680), .b(wfa_cout_681), .cin(wfa_s_682), .s(wfa_s_788), 
       .cout(wfa_cout_788));   // mult.v(3887)
    fa fa_789 (.a(wfa_cout_682), .b(wfa_cout_683), .cin(wfa_s_684), .s(wfa_s_789), 
       .cout(wfa_cout_789));   // mult.v(3888)
    fa fa_790 (.a(wfa_cout_684), .b(wfa_cout_685), .cin(wfa_s_686), .s(wfa_s_790), 
       .cout(wfa_cout_790));   // mult.v(3889)
    fa fa_791 (.a(wfa_cout_686), .b(wfa_cout_687), .cin(wfa_s_688), .s(wfa_s_791), 
       .cout(wfa_cout_791));   // mult.v(3890)
    fa fa_792 (.a(wfa_cout_688), .b(wfa_cout_689), .cin(wfa_s_690), .s(wfa_s_792), 
       .cout(wfa_cout_792));   // mult.v(3891)
    fa fa_793 (.a(wfa_cout_690), .b(wfa_cout_691), .cin(wfa_s_692), .s(wfa_s_793), 
       .cout(wfa_cout_793));   // mult.v(3892)
    fa fa_794 (.a(wfa_cout_692), .b(wfa_cout_693), .cin(wfa_s_694), .s(wfa_s_794), 
       .cout(wfa_cout_794));   // mult.v(3893)
    fa fa_795 (.a(wfa_cout_694), .b(wfa_cout_695), .cin(wfa_s_696), .s(wfa_s_795), 
       .cout(wfa_cout_795));   // mult.v(3894)
    fa fa_796 (.a(wfa_cout_696), .b(wfa_cout_697), .cin(wfa_s_698), .s(wfa_s_796), 
       .cout(wfa_cout_796));   // mult.v(3895)
    fa fa_797 (.a(wfa_cout_698), .b(wfa_cout_699), .cin(wfa_s_700), .s(wfa_s_797), 
       .cout(wfa_cout_797));   // mult.v(3896)
    fa fa_798 (.a(wfa_cout_700), .b(wfa_cout_701), .cin(wfa_s_702), .s(wfa_s_798), 
       .cout(wfa_cout_798));   // mult.v(3897)
    fa fa_799 (.a(wfa_cout_702), .b(wfa_cout_703), .cin(wfa_s_704), .s(wfa_s_799), 
       .cout(wfa_cout_799));   // mult.v(3898)
    fa fa_800 (.a(wfa_cout_704), .b(wfa_cout_705), .cin(wfa_s_706), .s(wfa_s_800), 
       .cout(wfa_cout_800));   // mult.v(3899)
    fa fa_801 (.a(wfa_cout_706), .b(wfa_cout_707), .cin(wfa_s_708), .s(wfa_s_801), 
       .cout(wfa_cout_801));   // mult.v(3900)
    fa fa_802 (.a(wfa_cout_708), .b(wfa_cout_709), .cin(wfa_s_710), .s(wfa_s_802), 
       .cout(wfa_cout_802));   // mult.v(3901)
    fa fa_803 (.a(wfa_cout_710), .b(wfa_cout_711), .cin(wfa_s_712), .s(wfa_s_803), 
       .cout(wfa_cout_803));   // mult.v(3902)
    fa fa_804 (.a(wfa_cout_712), .b(wfa_cout_713), .cin(wfa_s_714), .s(wfa_s_804), 
       .cout(wfa_cout_804));   // mult.v(3903)
    fa fa_805 (.a(wfa_cout_714), .b(wfa_cout_715), .cin(wfa_s_716), .s(wfa_s_805), 
       .cout(wfa_cout_805));   // mult.v(3904)
    fa fa_806 (.a(wfa_cout_716), .b(wfa_cout_717), .cin(wfa_s_718), .s(wfa_s_806), 
       .cout(wfa_cout_806));   // mult.v(3905)
    fa fa_807 (.a(wfa_cout_718), .b(wfa_cout_719), .cin(wfa_s_720), .s(wfa_s_807), 
       .cout(wfa_cout_807));   // mult.v(3906)
    fa fa_808 (.a(wfa_cout_720), .b(wfa_cout_721), .cin(wfa_s_722), .s(wfa_s_808), 
       .cout(wfa_cout_808));   // mult.v(3907)
    fa fa_809 (.a(wfa_cout_722), .b(wfa_cout_723), .cin(wfa_s_724), .s(wfa_s_809), 
       .cout(wfa_cout_809));   // mult.v(3908)
    fa fa_810 (.a(wfa_cout_724), .b(wfa_cout_725), .cin(wfa_s_726), .s(wfa_s_810), 
       .cout(wfa_cout_810));   // mult.v(3909)
    fa fa_811 (.a(wfa_cout_726), .b(wfa_cout_727), .cin(wfa_s_728), .s(wfa_s_811), 
       .cout(wfa_cout_811));   // mult.v(3910)
    fa fa_812 (.a(wfa_cout_728), .b(wfa_cout_729), .cin(wfa_s_730), .s(wfa_s_812), 
       .cout(wfa_cout_812));   // mult.v(3911)
    fa fa_813 (.a(wfa_cout_730), .b(wfa_cout_731), .cin(wfa_s_732), .s(wfa_s_813), 
       .cout(wfa_cout_813));   // mult.v(3912)
    fa fa_814 (.a(wfa_cout_732), .b(wfa_cout_733), .cin(wfa_s_734), .s(wfa_s_814), 
       .cout(wfa_cout_814));   // mult.v(3913)
    fa fa_815 (.a(wfa_cout_734), .b(wfa_cout_735), .cin(wfa_s_736), .s(wfa_s_815), 
       .cout(wfa_cout_815));   // mult.v(3914)
    fa fa_816 (.a(wfa_cout_736), .b(wfa_cout_737), .cin(wfa_s_738), .s(wfa_s_816), 
       .cout(wfa_cout_816));   // mult.v(3915)
    fa fa_817 (.a(wfa_cout_738), .b(wfa_cout_739), .cin(wfa_s_740), .s(wfa_s_817), 
       .cout(wfa_cout_817));   // mult.v(3916)
    fa fa_818 (.a(wfa_cout_740), .b(wfa_cout_741), .cin(wfa_s_742), .s(wfa_s_818), 
       .cout(wfa_cout_818));   // mult.v(3917)
    fa fa_819 (.a(wfa_cout_742), .b(wfa_cout_743), .cin(wfa_s_744), .s(wfa_s_819), 
       .cout(wfa_cout_819));   // mult.v(3918)
    fa fa_820 (.a(wfa_cout_744), .b(wfa_cout_745), .cin(wfa_s_746), .s(wfa_s_820), 
       .cout(wfa_cout_820));   // mult.v(3919)
    fa fa_821 (.a(wfa_cout_746), .b(wfa_cout_747), .cin(wfa_s_748), .s(wfa_s_821), 
       .cout(wfa_cout_821));   // mult.v(3920)
    fa fa_822 (.a(wfa_cout_748), .b(wfa_cout_749), .cin(wfa_s_750), .s(wfa_s_822), 
       .cout(wfa_cout_822));   // mult.v(3921)
    fa fa_823 (.a(wfa_cout_750), .b(wfa_cout_751), .cin(wfa_s_752), .s(wfa_s_823), 
       .cout(wfa_cout_823));   // mult.v(3922)
    fa fa_824 (.a(wfa_cout_752), .b(wfa_cout_753), .cin(wfa_s_754), .s(wfa_s_824), 
       .cout(wfa_cout_824));   // mult.v(3923)
    fa fa_825 (.a(wfa_cout_754), .b(wfa_cout_755), .cin(wfa_s_756), .s(wfa_s_825), 
       .cout(wfa_cout_825));   // mult.v(3924)
    fa fa_826 (.a(wfa_cout_756), .b(wfa_cout_757), .cin(wfa_s_758), .s(wfa_s_826), 
       .cout(wfa_cout_826));   // mult.v(3925)
    fa fa_827 (.a(wfa_cout_758), .b(wfa_cout_759), .cin(wfa_s_760), .s(wfa_s_827), 
       .cout(wfa_cout_827));   // mult.v(3926)
    fa fa_828 (.a(wfa_cout_760), .b(wfa_cout_761), .cin(wfa_s_762), .s(wfa_s_828), 
       .cout(wfa_cout_828));   // mult.v(3927)
    fa fa_829 (.a(wfa_cout_762), .b(wfa_cout_763), .cin(wfa_s_764), .s(wfa_s_829), 
       .cout(wfa_cout_829));   // mult.v(3928)
    fa fa_830 (.a(wfa_cout_764), .b(wfa_cout_765), .cin(wfa_s_766), .s(wfa_s_830), 
       .cout(wfa_cout_830));   // mult.v(3929)
    fa fa_831 (.a(wfa_cout_766), .b(wfa_cout_767), .cin(wfa_s_768), .s(wfa_s_831), 
       .cout(wfa_cout_831));   // mult.v(3930)
    fa fa_832 (.a(wfa_cout_768), .b(wfa_cout_769), .cin(wfa_s_770), .s(wfa_s_832), 
       .cout(wfa_cout_832));   // mult.v(3931)
    fa fa_833 (.a(wfa_cout_770), .b(wfa_cout_771), .cin(wfa_s_772), .s(wfa_s_833), 
       .cout(wfa_cout_833));   // mult.v(3932)
    fa fa_834 (.a(wfa_cout_772), .b(wfa_cout_773), .cin(wfa_s_774), .s(wfa_s_834), 
       .cout(wfa_cout_834));   // mult.v(3933)
    fa fa_835 (.a(wfa_cout_774), .b(wfa_cout_775), .cin(wfa_s_776), .s(wfa_s_835), 
       .cout(wfa_cout_835));   // mult.v(3934)
    fa fa_836 (.a(wfa_cout_776), .b(wfa_cout_777), .cin(wfa_s_778), .s(wfa_s_836), 
       .cout(wfa_cout_836));   // mult.v(3935)
    fa fa_837 (.a(wfa_cout_778), .b(wfa_cout_779), .cin(wfa_s_780), .s(wfa_s_837), 
       .cout(wfa_cout_837));   // mult.v(3936)
    and (wand_1020, a[31], b[28]) ;   // mult.v(3937)
    fa fa_838 (.a(wand_1020), .b(wfa_cout_780), .cin(wfa_cout_781), .s(wfa_s_838), 
       .cout(wfa_cout_838));   // mult.v(3938)
    and (wand_959, a[29], b[31]) ;   // mult.v(3939)
    and (wand_990, a[30], b[30]) ;   // mult.v(3940)
    and (wand_1021, a[31], b[29]) ;   // mult.v(3941)
    fa fa_839 (.a(wand_959), .b(wand_990), .cin(wand_1021), .s(wfa_s_839), 
       .cout(wfa_cout_839));   // mult.v(3942)
    and (wand_2, a[0], b[2]) ;   // mult.v(3943)
    and (wand_33, a[1], b[1]) ;   // mult.v(3944)
    ha ha_30 (.a(wand_2), .b(wand_33), .s(wha_s_30), .c(wha_c_30));   // mult.v(3945)
    and (wand_65, a[2], b[1]) ;   // mult.v(3946)
    and (wand_96, a[3], b[0]) ;   // mult.v(3947)
    fa fa_840 (.a(wand_65), .b(wand_96), .cin(wha_s_29), .s(wfa_s_840), 
       .cout(wfa_cout_840));   // mult.v(3948)
    fa fa_841 (.a(wha_s_27), .b(wha_c_29), .cin(wfa_s_783), .s(wfa_s_841), 
       .cout(wfa_cout_841));   // mult.v(3949)
    fa fa_842 (.a(wha_s_28), .b(wfa_cout_783), .cin(wfa_s_784), .s(wfa_s_842), 
       .cout(wfa_cout_842));   // mult.v(3950)
    fa fa_843 (.a(wfa_s_677), .b(wfa_cout_784), .cin(wfa_s_785), .s(wfa_s_843), 
       .cout(wfa_cout_843));   // mult.v(3951)
    fa fa_844 (.a(wfa_s_679), .b(wfa_cout_785), .cin(wfa_s_786), .s(wfa_s_844), 
       .cout(wfa_cout_844));   // mult.v(3952)
    fa fa_845 (.a(wfa_s_681), .b(wfa_cout_786), .cin(wfa_s_787), .s(wfa_s_845), 
       .cout(wfa_cout_845));   // mult.v(3953)
    fa fa_846 (.a(wfa_s_683), .b(wfa_cout_787), .cin(wfa_s_788), .s(wfa_s_846), 
       .cout(wfa_cout_846));   // mult.v(3954)
    fa fa_847 (.a(wfa_s_685), .b(wfa_cout_788), .cin(wfa_s_789), .s(wfa_s_847), 
       .cout(wfa_cout_847));   // mult.v(3955)
    fa fa_848 (.a(wfa_s_687), .b(wfa_cout_789), .cin(wfa_s_790), .s(wfa_s_848), 
       .cout(wfa_cout_848));   // mult.v(3956)
    fa fa_849 (.a(wfa_s_689), .b(wfa_cout_790), .cin(wfa_s_791), .s(wfa_s_849), 
       .cout(wfa_cout_849));   // mult.v(3957)
    fa fa_850 (.a(wfa_s_691), .b(wfa_cout_791), .cin(wfa_s_792), .s(wfa_s_850), 
       .cout(wfa_cout_850));   // mult.v(3958)
    fa fa_851 (.a(wfa_s_693), .b(wfa_cout_792), .cin(wfa_s_793), .s(wfa_s_851), 
       .cout(wfa_cout_851));   // mult.v(3959)
    fa fa_852 (.a(wfa_s_695), .b(wfa_cout_793), .cin(wfa_s_794), .s(wfa_s_852), 
       .cout(wfa_cout_852));   // mult.v(3960)
    fa fa_853 (.a(wfa_s_697), .b(wfa_cout_794), .cin(wfa_s_795), .s(wfa_s_853), 
       .cout(wfa_cout_853));   // mult.v(3961)
    fa fa_854 (.a(wfa_s_699), .b(wfa_cout_795), .cin(wfa_s_796), .s(wfa_s_854), 
       .cout(wfa_cout_854));   // mult.v(3962)
    fa fa_855 (.a(wfa_s_701), .b(wfa_cout_796), .cin(wfa_s_797), .s(wfa_s_855), 
       .cout(wfa_cout_855));   // mult.v(3963)
    fa fa_856 (.a(wfa_s_703), .b(wfa_cout_797), .cin(wfa_s_798), .s(wfa_s_856), 
       .cout(wfa_cout_856));   // mult.v(3964)
    fa fa_857 (.a(wfa_s_705), .b(wfa_cout_798), .cin(wfa_s_799), .s(wfa_s_857), 
       .cout(wfa_cout_857));   // mult.v(3965)
    fa fa_858 (.a(wfa_s_707), .b(wfa_cout_799), .cin(wfa_s_800), .s(wfa_s_858), 
       .cout(wfa_cout_858));   // mult.v(3966)
    fa fa_859 (.a(wfa_s_709), .b(wfa_cout_800), .cin(wfa_s_801), .s(wfa_s_859), 
       .cout(wfa_cout_859));   // mult.v(3967)
    fa fa_860 (.a(wfa_s_711), .b(wfa_cout_801), .cin(wfa_s_802), .s(wfa_s_860), 
       .cout(wfa_cout_860));   // mult.v(3968)
    fa fa_861 (.a(wfa_s_713), .b(wfa_cout_802), .cin(wfa_s_803), .s(wfa_s_861), 
       .cout(wfa_cout_861));   // mult.v(3969)
    fa fa_862 (.a(wfa_s_715), .b(wfa_cout_803), .cin(wfa_s_804), .s(wfa_s_862), 
       .cout(wfa_cout_862));   // mult.v(3970)
    fa fa_863 (.a(wfa_s_717), .b(wfa_cout_804), .cin(wfa_s_805), .s(wfa_s_863), 
       .cout(wfa_cout_863));   // mult.v(3971)
    fa fa_864 (.a(wfa_s_719), .b(wfa_cout_805), .cin(wfa_s_806), .s(wfa_s_864), 
       .cout(wfa_cout_864));   // mult.v(3972)
    fa fa_865 (.a(wfa_s_721), .b(wfa_cout_806), .cin(wfa_s_807), .s(wfa_s_865), 
       .cout(wfa_cout_865));   // mult.v(3973)
    fa fa_866 (.a(wfa_s_723), .b(wfa_cout_807), .cin(wfa_s_808), .s(wfa_s_866), 
       .cout(wfa_cout_866));   // mult.v(3974)
    fa fa_867 (.a(wfa_s_725), .b(wfa_cout_808), .cin(wfa_s_809), .s(wfa_s_867), 
       .cout(wfa_cout_867));   // mult.v(3975)
    fa fa_868 (.a(wfa_s_727), .b(wfa_cout_809), .cin(wfa_s_810), .s(wfa_s_868), 
       .cout(wfa_cout_868));   // mult.v(3976)
    fa fa_869 (.a(wfa_s_729), .b(wfa_cout_810), .cin(wfa_s_811), .s(wfa_s_869), 
       .cout(wfa_cout_869));   // mult.v(3977)
    fa fa_870 (.a(wfa_s_731), .b(wfa_cout_811), .cin(wfa_s_812), .s(wfa_s_870), 
       .cout(wfa_cout_870));   // mult.v(3978)
    fa fa_871 (.a(wfa_s_733), .b(wfa_cout_812), .cin(wfa_s_813), .s(wfa_s_871), 
       .cout(wfa_cout_871));   // mult.v(3979)
    fa fa_872 (.a(wfa_s_735), .b(wfa_cout_813), .cin(wfa_s_814), .s(wfa_s_872), 
       .cout(wfa_cout_872));   // mult.v(3980)
    fa fa_873 (.a(wfa_s_737), .b(wfa_cout_814), .cin(wfa_s_815), .s(wfa_s_873), 
       .cout(wfa_cout_873));   // mult.v(3981)
    fa fa_874 (.a(wfa_s_739), .b(wfa_cout_815), .cin(wfa_s_816), .s(wfa_s_874), 
       .cout(wfa_cout_874));   // mult.v(3982)
    fa fa_875 (.a(wfa_s_741), .b(wfa_cout_816), .cin(wfa_s_817), .s(wfa_s_875), 
       .cout(wfa_cout_875));   // mult.v(3983)
    fa fa_876 (.a(wfa_s_743), .b(wfa_cout_817), .cin(wfa_s_818), .s(wfa_s_876), 
       .cout(wfa_cout_876));   // mult.v(3984)
    fa fa_877 (.a(wfa_s_745), .b(wfa_cout_818), .cin(wfa_s_819), .s(wfa_s_877), 
       .cout(wfa_cout_877));   // mult.v(3985)
    fa fa_878 (.a(wfa_s_747), .b(wfa_cout_819), .cin(wfa_s_820), .s(wfa_s_878), 
       .cout(wfa_cout_878));   // mult.v(3986)
    fa fa_879 (.a(wfa_s_749), .b(wfa_cout_820), .cin(wfa_s_821), .s(wfa_s_879), 
       .cout(wfa_cout_879));   // mult.v(3987)
    fa fa_880 (.a(wfa_s_751), .b(wfa_cout_821), .cin(wfa_s_822), .s(wfa_s_880), 
       .cout(wfa_cout_880));   // mult.v(3988)
    fa fa_881 (.a(wfa_s_753), .b(wfa_cout_822), .cin(wfa_s_823), .s(wfa_s_881), 
       .cout(wfa_cout_881));   // mult.v(3989)
    fa fa_882 (.a(wfa_s_755), .b(wfa_cout_823), .cin(wfa_s_824), .s(wfa_s_882), 
       .cout(wfa_cout_882));   // mult.v(3990)
    fa fa_883 (.a(wfa_s_757), .b(wfa_cout_824), .cin(wfa_s_825), .s(wfa_s_883), 
       .cout(wfa_cout_883));   // mult.v(3991)
    fa fa_884 (.a(wfa_s_759), .b(wfa_cout_825), .cin(wfa_s_826), .s(wfa_s_884), 
       .cout(wfa_cout_884));   // mult.v(3992)
    fa fa_885 (.a(wfa_s_761), .b(wfa_cout_826), .cin(wfa_s_827), .s(wfa_s_885), 
       .cout(wfa_cout_885));   // mult.v(3993)
    fa fa_886 (.a(wfa_s_763), .b(wfa_cout_827), .cin(wfa_s_828), .s(wfa_s_886), 
       .cout(wfa_cout_886));   // mult.v(3994)
    fa fa_887 (.a(wfa_s_765), .b(wfa_cout_828), .cin(wfa_s_829), .s(wfa_s_887), 
       .cout(wfa_cout_887));   // mult.v(3995)
    fa fa_888 (.a(wfa_s_767), .b(wfa_cout_829), .cin(wfa_s_830), .s(wfa_s_888), 
       .cout(wfa_cout_888));   // mult.v(3996)
    fa fa_889 (.a(wfa_s_769), .b(wfa_cout_830), .cin(wfa_s_831), .s(wfa_s_889), 
       .cout(wfa_cout_889));   // mult.v(3997)
    fa fa_890 (.a(wfa_s_771), .b(wfa_cout_831), .cin(wfa_s_832), .s(wfa_s_890), 
       .cout(wfa_cout_890));   // mult.v(3998)
    fa fa_891 (.a(wfa_s_773), .b(wfa_cout_832), .cin(wfa_s_833), .s(wfa_s_891), 
       .cout(wfa_cout_891));   // mult.v(3999)
    fa fa_892 (.a(wfa_s_775), .b(wfa_cout_833), .cin(wfa_s_834), .s(wfa_s_892), 
       .cout(wfa_cout_892));   // mult.v(4000)
    fa fa_893 (.a(wfa_s_777), .b(wfa_cout_834), .cin(wfa_s_835), .s(wfa_s_893), 
       .cout(wfa_cout_893));   // mult.v(4001)
    fa fa_894 (.a(wfa_s_779), .b(wfa_cout_835), .cin(wfa_s_836), .s(wfa_s_894), 
       .cout(wfa_cout_894));   // mult.v(4002)
    fa fa_895 (.a(wfa_s_781), .b(wfa_cout_836), .cin(wfa_s_837), .s(wfa_s_895), 
       .cout(wfa_cout_895));   // mult.v(4003)
    fa fa_896 (.a(wfa_s_782), .b(wfa_cout_837), .cin(wfa_s_838), .s(wfa_s_896), 
       .cout(wfa_cout_896));   // mult.v(4004)
    fa fa_897 (.a(wfa_cout_782), .b(wfa_cout_838), .cin(wfa_s_839), .s(wfa_s_897), 
       .cout(wfa_cout_897));   // mult.v(4005)
    and (wand_991, a[30], b[31]) ;   // mult.v(4006)
    and (wand_1022, a[31], b[30]) ;   // mult.v(4007)
    fa fa_898 (.a(wand_991), .b(wand_1022), .cin(wfa_cout_839), .s(wfa_s_898), 
       .cout(wfa_cout_898));   // mult.v(4008)
    and (wand_1, a[0], b[1]) ;   // mult.v(4009)
    and (wand_32, a[1], b[0]) ;   // mult.v(4010)
    ha ha_31 (.a(wand_1), .b(wand_32), .s(m[1]), .c(wha_c_31));   // mult.v(4011)
    and (wand_64, a[2], b[0]) ;   // mult.v(4012)
    fa fa_899 (.a(wand_64), .b(wha_s_30), .cin(wha_c_31), .s(m[2]), 
       .cout(wfa_cout_899));   // mult.v(4013)
    fa fa_900 (.a(wha_c_30), .b(wfa_s_840), .cin(wfa_cout_899), .s(m[3]), 
       .cout(wfa_cout_900));   // mult.v(4014)
    fa fa_901 (.a(wfa_cout_840), .b(wfa_s_841), .cin(wfa_cout_900), .s(m[4]), 
       .cout(wfa_cout_901));   // mult.v(4015)
    fa fa_902 (.a(wfa_cout_841), .b(wfa_s_842), .cin(wfa_cout_901), .s(m[5]), 
       .cout(wfa_cout_902));   // mult.v(4016)
    fa fa_903 (.a(wfa_cout_842), .b(wfa_s_843), .cin(wfa_cout_902), .s(m[6]), 
       .cout(wfa_cout_903));   // mult.v(4017)
    fa fa_904 (.a(wfa_cout_843), .b(wfa_s_844), .cin(wfa_cout_903), .s(m[7]), 
       .cout(wfa_cout_904));   // mult.v(4018)
    fa fa_905 (.a(wfa_cout_844), .b(wfa_s_845), .cin(wfa_cout_904), .s(m[8]), 
       .cout(wfa_cout_905));   // mult.v(4019)
    fa fa_906 (.a(wfa_cout_845), .b(wfa_s_846), .cin(wfa_cout_905), .s(m[9]), 
       .cout(wfa_cout_906));   // mult.v(4020)
    fa fa_907 (.a(wfa_cout_846), .b(wfa_s_847), .cin(wfa_cout_906), .s(m[10]), 
       .cout(wfa_cout_907));   // mult.v(4021)
    fa fa_908 (.a(wfa_cout_847), .b(wfa_s_848), .cin(wfa_cout_907), .s(m[11]), 
       .cout(wfa_cout_908));   // mult.v(4022)
    fa fa_909 (.a(wfa_cout_848), .b(wfa_s_849), .cin(wfa_cout_908), .s(m[12]), 
       .cout(wfa_cout_909));   // mult.v(4023)
    fa fa_910 (.a(wfa_cout_849), .b(wfa_s_850), .cin(wfa_cout_909), .s(m[13]), 
       .cout(wfa_cout_910));   // mult.v(4024)
    fa fa_911 (.a(wfa_cout_850), .b(wfa_s_851), .cin(wfa_cout_910), .s(m[14]), 
       .cout(wfa_cout_911));   // mult.v(4025)
    fa fa_912 (.a(wfa_cout_851), .b(wfa_s_852), .cin(wfa_cout_911), .s(m[15]), 
       .cout(wfa_cout_912));   // mult.v(4026)
    fa fa_913 (.a(wfa_cout_852), .b(wfa_s_853), .cin(wfa_cout_912), .s(m[16]), 
       .cout(wfa_cout_913));   // mult.v(4027)
    fa fa_914 (.a(wfa_cout_853), .b(wfa_s_854), .cin(wfa_cout_913), .s(m[17]), 
       .cout(wfa_cout_914));   // mult.v(4028)
    fa fa_915 (.a(wfa_cout_854), .b(wfa_s_855), .cin(wfa_cout_914), .s(m[18]), 
       .cout(wfa_cout_915));   // mult.v(4029)
    fa fa_916 (.a(wfa_cout_855), .b(wfa_s_856), .cin(wfa_cout_915), .s(m[19]), 
       .cout(wfa_cout_916));   // mult.v(4030)
    fa fa_917 (.a(wfa_cout_856), .b(wfa_s_857), .cin(wfa_cout_916), .s(m[20]), 
       .cout(wfa_cout_917));   // mult.v(4031)
    fa fa_918 (.a(wfa_cout_857), .b(wfa_s_858), .cin(wfa_cout_917), .s(m[21]), 
       .cout(wfa_cout_918));   // mult.v(4032)
    fa fa_919 (.a(wfa_cout_858), .b(wfa_s_859), .cin(wfa_cout_918), .s(m[22]), 
       .cout(wfa_cout_919));   // mult.v(4033)
    fa fa_920 (.a(wfa_cout_859), .b(wfa_s_860), .cin(wfa_cout_919), .s(m[23]), 
       .cout(wfa_cout_920));   // mult.v(4034)
    fa fa_921 (.a(wfa_cout_860), .b(wfa_s_861), .cin(wfa_cout_920), .s(m[24]), 
       .cout(wfa_cout_921));   // mult.v(4035)
    fa fa_922 (.a(wfa_cout_861), .b(wfa_s_862), .cin(wfa_cout_921), .s(m[25]), 
       .cout(wfa_cout_922));   // mult.v(4036)
    fa fa_923 (.a(wfa_cout_862), .b(wfa_s_863), .cin(wfa_cout_922), .s(m[26]), 
       .cout(wfa_cout_923));   // mult.v(4037)
    fa fa_924 (.a(wfa_cout_863), .b(wfa_s_864), .cin(wfa_cout_923), .s(m[27]), 
       .cout(wfa_cout_924));   // mult.v(4038)
    fa fa_925 (.a(wfa_cout_864), .b(wfa_s_865), .cin(wfa_cout_924), .s(m[28]), 
       .cout(wfa_cout_925));   // mult.v(4039)
    fa fa_926 (.a(wfa_cout_865), .b(wfa_s_866), .cin(wfa_cout_925), .s(m[29]), 
       .cout(wfa_cout_926));   // mult.v(4040)
    fa fa_927 (.a(wfa_cout_866), .b(wfa_s_867), .cin(wfa_cout_926), .s(m[30]), 
       .cout(wfa_cout_927));   // mult.v(4041)
    fa fa_928 (.a(wfa_cout_867), .b(wfa_s_868), .cin(wfa_cout_927), .s(m[31]), 
       .cout(wfa_cout_928));   // mult.v(4042)
    fa fa_929 (.a(wfa_cout_868), .b(wfa_s_869), .cin(wfa_cout_928), .s(m[32]), 
       .cout(wfa_cout_929));   // mult.v(4043)
    fa fa_930 (.a(wfa_cout_869), .b(wfa_s_870), .cin(wfa_cout_929), .s(m[33]), 
       .cout(wfa_cout_930));   // mult.v(4044)
    fa fa_931 (.a(wfa_cout_870), .b(wfa_s_871), .cin(wfa_cout_930), .s(m[34]), 
       .cout(wfa_cout_931));   // mult.v(4045)
    fa fa_932 (.a(wfa_cout_871), .b(wfa_s_872), .cin(wfa_cout_931), .s(m[35]), 
       .cout(wfa_cout_932));   // mult.v(4046)
    fa fa_933 (.a(wfa_cout_872), .b(wfa_s_873), .cin(wfa_cout_932), .s(m[36]), 
       .cout(wfa_cout_933));   // mult.v(4047)
    fa fa_934 (.a(wfa_cout_873), .b(wfa_s_874), .cin(wfa_cout_933), .s(m[37]), 
       .cout(wfa_cout_934));   // mult.v(4048)
    fa fa_935 (.a(wfa_cout_874), .b(wfa_s_875), .cin(wfa_cout_934), .s(m[38]), 
       .cout(wfa_cout_935));   // mult.v(4049)
    fa fa_936 (.a(wfa_cout_875), .b(wfa_s_876), .cin(wfa_cout_935), .s(m[39]), 
       .cout(wfa_cout_936));   // mult.v(4050)
    fa fa_937 (.a(wfa_cout_876), .b(wfa_s_877), .cin(wfa_cout_936), .s(m[40]), 
       .cout(wfa_cout_937));   // mult.v(4051)
    fa fa_938 (.a(wfa_cout_877), .b(wfa_s_878), .cin(wfa_cout_937), .s(m[41]), 
       .cout(wfa_cout_938));   // mult.v(4052)
    fa fa_939 (.a(wfa_cout_878), .b(wfa_s_879), .cin(wfa_cout_938), .s(m[42]), 
       .cout(wfa_cout_939));   // mult.v(4053)
    fa fa_940 (.a(wfa_cout_879), .b(wfa_s_880), .cin(wfa_cout_939), .s(m[43]), 
       .cout(wfa_cout_940));   // mult.v(4054)
    fa fa_941 (.a(wfa_cout_880), .b(wfa_s_881), .cin(wfa_cout_940), .s(m[44]), 
       .cout(wfa_cout_941));   // mult.v(4055)
    fa fa_942 (.a(wfa_cout_881), .b(wfa_s_882), .cin(wfa_cout_941), .s(m[45]), 
       .cout(wfa_cout_942));   // mult.v(4056)
    fa fa_943 (.a(wfa_cout_882), .b(wfa_s_883), .cin(wfa_cout_942), .s(m[46]), 
       .cout(wfa_cout_943));   // mult.v(4057)
    fa fa_944 (.a(wfa_cout_883), .b(wfa_s_884), .cin(wfa_cout_943), .s(m[47]), 
       .cout(wfa_cout_944));   // mult.v(4058)
    fa fa_945 (.a(wfa_cout_884), .b(wfa_s_885), .cin(wfa_cout_944), .s(m[48]), 
       .cout(wfa_cout_945));   // mult.v(4059)
    fa fa_946 (.a(wfa_cout_885), .b(wfa_s_886), .cin(wfa_cout_945), .s(m[49]), 
       .cout(wfa_cout_946));   // mult.v(4060)
    fa fa_947 (.a(wfa_cout_886), .b(wfa_s_887), .cin(wfa_cout_946), .s(m[50]), 
       .cout(wfa_cout_947));   // mult.v(4061)
    fa fa_948 (.a(wfa_cout_887), .b(wfa_s_888), .cin(wfa_cout_947), .s(m[51]), 
       .cout(wfa_cout_948));   // mult.v(4062)
    fa fa_949 (.a(wfa_cout_888), .b(wfa_s_889), .cin(wfa_cout_948), .s(m[52]), 
       .cout(wfa_cout_949));   // mult.v(4063)
    fa fa_950 (.a(wfa_cout_889), .b(wfa_s_890), .cin(wfa_cout_949), .s(m[53]), 
       .cout(wfa_cout_950));   // mult.v(4064)
    fa fa_951 (.a(wfa_cout_890), .b(wfa_s_891), .cin(wfa_cout_950), .s(m[54]), 
       .cout(wfa_cout_951));   // mult.v(4065)
    fa fa_952 (.a(wfa_cout_891), .b(wfa_s_892), .cin(wfa_cout_951), .s(m[55]), 
       .cout(wfa_cout_952));   // mult.v(4066)
    fa fa_953 (.a(wfa_cout_892), .b(wfa_s_893), .cin(wfa_cout_952), .s(m[56]), 
       .cout(wfa_cout_953));   // mult.v(4067)
    fa fa_954 (.a(wfa_cout_893), .b(wfa_s_894), .cin(wfa_cout_953), .s(m[57]), 
       .cout(wfa_cout_954));   // mult.v(4068)
    fa fa_955 (.a(wfa_cout_894), .b(wfa_s_895), .cin(wfa_cout_954), .s(m[58]), 
       .cout(wfa_cout_955));   // mult.v(4069)
    fa fa_956 (.a(wfa_cout_895), .b(wfa_s_896), .cin(wfa_cout_955), .s(m[59]), 
       .cout(wfa_cout_956));   // mult.v(4070)
    fa fa_957 (.a(wfa_cout_896), .b(wfa_s_897), .cin(wfa_cout_956), .s(m[60]), 
       .cout(wfa_cout_957));   // mult.v(4071)
    fa fa_958 (.a(wfa_cout_897), .b(wfa_s_898), .cin(wfa_cout_957), .s(m[61]), 
       .cout(wfa_cout_958));   // mult.v(4072)
    and (wand_1023, a[31], b[31]) ;   // mult.v(4073)
    fa fa_959 (.a(wand_1023), .b(wfa_cout_898), .cin(wfa_cout_958), .s(m[62]), 
       .cout(m[63]));   // mult.v(4074)
    and (m[0], a[0], b[0]) ;   // mult.v(4075)
    
endmodule

//
// Verific Verilog Description of module ha
//

module ha (a, b, s, c);   // mult.v(25)
    input a;   // mult.v(26)
    input b;   // mult.v(27)
    output s;   // mult.v(29)
    output c;   // mult.v(30)
    
    
    xor (s, a, b) ;   // mult.v(32)
    and (c, a, b) ;   // mult.v(33)
    
endmodule

//
// Verific Verilog Description of module fa
//

module fa (a, b, cin, s, cout);   // mult.v(7)
    input a;   // mult.v(8)
    input b;   // mult.v(9)
    input cin;   // mult.v(10)
    output s;   // mult.v(12)
    output cout;   // mult.v(13)
    
    wire w1;   // mult.v(15)
    wire w2;   // mult.v(15)
    wire w3;   // mult.v(15)
    
    xor (w1, a, b) ;   // mult.v(17)
    xor (s, w1, cin) ;   // mult.v(18)
    and (w2, a, b) ;   // mult.v(20)
    and (w3, w1, cin) ;   // mult.v(21)
    or (cout, w2, w3) ;   // mult.v(22)
    
endmodule

//
// Verific Verilog Description of module bitwise_32
//

module bitwise_32 (q, z, a, b, op);   // alu.v(39)
    output [31:0]q;   // alu.v(43)
    output z;   // alu.v(44)
    input [31:0]a;   // alu.v(40)
    input [31:0]b;   // alu.v(40)
    input [2:0]op;   // alu.v(41)
    
    
    wire n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
        n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, 
        n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, 
        n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
        n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, 
        n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, 
        n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, 
        n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, 
        n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
        n96, n97, n98, n99, n100, n101, n102, n103, n104, 
        n105, n106, n107, n108, n109, n110, n111, n112, n113, 
        n114, n115, n116, n117, n118, n119, n120, n121, n122, 
        n123, n124, n125, n126, n127, n128, n129, n130, n131, 
        n132, n165, n166, n167, n168, n169, n170, n171, n172, 
        n173, n174, n175, n176, n177, n178, n179, n180, n181, 
        n182, n183, n184, n185, n186, n187, n188, n189, n190, 
        n191, n192, n193, n194, n195, n196, n229, n230, n231, 
        n232, n233, n234, n235, n236, n237, n238, n239, n240, 
        n241, n242, n243, n244, n245, n246, n247, n248, n249, 
        n250, n251, n252, n253, n254, n255, n256, n257, n258, 
        n259, n260, n293, n294, n295, n296, n297, n298, n299, 
        n300, n301, n302, n303, n304, n305, n306, n307, n308, 
        n309, n310, n311, n312, n313, n314, n315, n316, n317, 
        n318, n319, n320, n321, n322, n323, n324, n325, n326, 
        n327, n328, n329, n330, n331, n332, n333, n334, n335, 
        n336, n337, n338, n339, n340, n341, n342, n343, n344, 
        n345, n346, n347, n348, n349, n350, n351, n352, n353, 
        n354, n355, n356;
    
    nor (z, q[31], q[30], q[29], q[28], q[27], q[26], q[25], 
        q[24], q[23], q[22], q[21], q[20], q[19], q[18], q[17], 
        q[16], q[15], q[14], q[13], q[12], q[11], q[10], q[9], 
        q[8], q[7], q[6], q[5], q[4], q[3], q[2], q[1], q[0]) ;   // alu.v(46)
    not (n5, a[31]) ;   // alu.v(50)
    not (n6, a[30]) ;   // alu.v(50)
    not (n7, a[29]) ;   // alu.v(50)
    not (n8, a[28]) ;   // alu.v(50)
    not (n9, a[27]) ;   // alu.v(50)
    not (n10, a[26]) ;   // alu.v(50)
    not (n11, a[25]) ;   // alu.v(50)
    not (n12, a[24]) ;   // alu.v(50)
    not (n13, a[23]) ;   // alu.v(50)
    not (n14, a[22]) ;   // alu.v(50)
    not (n15, a[21]) ;   // alu.v(50)
    not (n16, a[20]) ;   // alu.v(50)
    not (n17, a[19]) ;   // alu.v(50)
    not (n18, a[18]) ;   // alu.v(50)
    not (n19, a[17]) ;   // alu.v(50)
    not (n20, a[16]) ;   // alu.v(50)
    not (n21, a[15]) ;   // alu.v(50)
    not (n22, a[14]) ;   // alu.v(50)
    not (n23, a[13]) ;   // alu.v(50)
    not (n24, a[12]) ;   // alu.v(50)
    not (n25, a[11]) ;   // alu.v(50)
    not (n26, a[10]) ;   // alu.v(50)
    not (n27, a[9]) ;   // alu.v(50)
    not (n28, a[8]) ;   // alu.v(50)
    not (n29, a[7]) ;   // alu.v(50)
    not (n30, a[6]) ;   // alu.v(50)
    not (n31, a[5]) ;   // alu.v(50)
    not (n32, a[4]) ;   // alu.v(50)
    not (n33, a[3]) ;   // alu.v(50)
    not (n34, a[2]) ;   // alu.v(50)
    not (n35, a[1]) ;   // alu.v(50)
    not (n36, a[0]) ;   // alu.v(50)
    and (n37, a[0], b[0]) ;   // alu.v(51)
    and (n38, a[1], b[1]) ;   // alu.v(51)
    and (n39, a[2], b[2]) ;   // alu.v(51)
    and (n40, a[3], b[3]) ;   // alu.v(51)
    and (n41, a[4], b[4]) ;   // alu.v(51)
    and (n42, a[5], b[5]) ;   // alu.v(51)
    and (n43, a[6], b[6]) ;   // alu.v(51)
    and (n44, a[7], b[7]) ;   // alu.v(51)
    and (n45, a[8], b[8]) ;   // alu.v(51)
    and (n46, a[9], b[9]) ;   // alu.v(51)
    and (n47, a[10], b[10]) ;   // alu.v(51)
    and (n48, a[11], b[11]) ;   // alu.v(51)
    and (n49, a[12], b[12]) ;   // alu.v(51)
    and (n50, a[13], b[13]) ;   // alu.v(51)
    and (n51, a[14], b[14]) ;   // alu.v(51)
    and (n52, a[15], b[15]) ;   // alu.v(51)
    and (n53, a[16], b[16]) ;   // alu.v(51)
    and (n54, a[17], b[17]) ;   // alu.v(51)
    and (n55, a[18], b[18]) ;   // alu.v(51)
    and (n56, a[19], b[19]) ;   // alu.v(51)
    and (n57, a[20], b[20]) ;   // alu.v(51)
    and (n58, a[21], b[21]) ;   // alu.v(51)
    and (n59, a[22], b[22]) ;   // alu.v(51)
    and (n60, a[23], b[23]) ;   // alu.v(51)
    and (n61, a[24], b[24]) ;   // alu.v(51)
    and (n62, a[25], b[25]) ;   // alu.v(51)
    and (n63, a[26], b[26]) ;   // alu.v(51)
    and (n64, a[27], b[27]) ;   // alu.v(51)
    and (n65, a[28], b[28]) ;   // alu.v(51)
    and (n66, a[29], b[29]) ;   // alu.v(51)
    and (n67, a[30], b[30]) ;   // alu.v(51)
    and (n68, a[31], b[31]) ;   // alu.v(51)
    or (n69, a[0], b[0]) ;   // alu.v(52)
    or (n70, a[1], b[1]) ;   // alu.v(52)
    or (n71, a[2], b[2]) ;   // alu.v(52)
    or (n72, a[3], b[3]) ;   // alu.v(52)
    or (n73, a[4], b[4]) ;   // alu.v(52)
    or (n74, a[5], b[5]) ;   // alu.v(52)
    or (n75, a[6], b[6]) ;   // alu.v(52)
    or (n76, a[7], b[7]) ;   // alu.v(52)
    or (n77, a[8], b[8]) ;   // alu.v(52)
    or (n78, a[9], b[9]) ;   // alu.v(52)
    or (n79, a[10], b[10]) ;   // alu.v(52)
    or (n80, a[11], b[11]) ;   // alu.v(52)
    or (n81, a[12], b[12]) ;   // alu.v(52)
    or (n82, a[13], b[13]) ;   // alu.v(52)
    or (n83, a[14], b[14]) ;   // alu.v(52)
    or (n84, a[15], b[15]) ;   // alu.v(52)
    or (n85, a[16], b[16]) ;   // alu.v(52)
    or (n86, a[17], b[17]) ;   // alu.v(52)
    or (n87, a[18], b[18]) ;   // alu.v(52)
    or (n88, a[19], b[19]) ;   // alu.v(52)
    or (n89, a[20], b[20]) ;   // alu.v(52)
    or (n90, a[21], b[21]) ;   // alu.v(52)
    or (n91, a[22], b[22]) ;   // alu.v(52)
    or (n92, a[23], b[23]) ;   // alu.v(52)
    or (n93, a[24], b[24]) ;   // alu.v(52)
    or (n94, a[25], b[25]) ;   // alu.v(52)
    or (n95, a[26], b[26]) ;   // alu.v(52)
    or (n96, a[27], b[27]) ;   // alu.v(52)
    or (n97, a[28], b[28]) ;   // alu.v(52)
    or (n98, a[29], b[29]) ;   // alu.v(52)
    or (n99, a[30], b[30]) ;   // alu.v(52)
    or (n100, a[31], b[31]) ;   // alu.v(52)
    xor (n101, a[0], b[0]) ;   // alu.v(53)
    xor (n102, a[1], b[1]) ;   // alu.v(53)
    xor (n103, a[2], b[2]) ;   // alu.v(53)
    xor (n104, a[3], b[3]) ;   // alu.v(53)
    xor (n105, a[4], b[4]) ;   // alu.v(53)
    xor (n106, a[5], b[5]) ;   // alu.v(53)
    xor (n107, a[6], b[6]) ;   // alu.v(53)
    xor (n108, a[7], b[7]) ;   // alu.v(53)
    xor (n109, a[8], b[8]) ;   // alu.v(53)
    xor (n110, a[9], b[9]) ;   // alu.v(53)
    xor (n111, a[10], b[10]) ;   // alu.v(53)
    xor (n112, a[11], b[11]) ;   // alu.v(53)
    xor (n113, a[12], b[12]) ;   // alu.v(53)
    xor (n114, a[13], b[13]) ;   // alu.v(53)
    xor (n115, a[14], b[14]) ;   // alu.v(53)
    xor (n116, a[15], b[15]) ;   // alu.v(53)
    xor (n117, a[16], b[16]) ;   // alu.v(53)
    xor (n118, a[17], b[17]) ;   // alu.v(53)
    xor (n119, a[18], b[18]) ;   // alu.v(53)
    xor (n120, a[19], b[19]) ;   // alu.v(53)
    xor (n121, a[20], b[20]) ;   // alu.v(53)
    xor (n122, a[21], b[21]) ;   // alu.v(53)
    xor (n123, a[22], b[22]) ;   // alu.v(53)
    xor (n124, a[23], b[23]) ;   // alu.v(53)
    xor (n125, a[24], b[24]) ;   // alu.v(53)
    xor (n126, a[25], b[25]) ;   // alu.v(53)
    xor (n127, a[26], b[26]) ;   // alu.v(53)
    xor (n128, a[27], b[27]) ;   // alu.v(53)
    xor (n129, a[28], b[28]) ;   // alu.v(53)
    xor (n130, a[29], b[29]) ;   // alu.v(53)
    xor (n131, a[30], b[30]) ;   // alu.v(53)
    xor (n132, a[31], b[31]) ;   // alu.v(53)
    not (n165, n68) ;   // alu.v(54)
    not (n166, n67) ;   // alu.v(54)
    not (n167, n66) ;   // alu.v(54)
    not (n168, n65) ;   // alu.v(54)
    not (n169, n64) ;   // alu.v(54)
    not (n170, n63) ;   // alu.v(54)
    not (n171, n62) ;   // alu.v(54)
    not (n172, n61) ;   // alu.v(54)
    not (n173, n60) ;   // alu.v(54)
    not (n174, n59) ;   // alu.v(54)
    not (n175, n58) ;   // alu.v(54)
    not (n176, n57) ;   // alu.v(54)
    not (n177, n56) ;   // alu.v(54)
    not (n178, n55) ;   // alu.v(54)
    not (n179, n54) ;   // alu.v(54)
    not (n180, n53) ;   // alu.v(54)
    not (n181, n52) ;   // alu.v(54)
    not (n182, n51) ;   // alu.v(54)
    not (n183, n50) ;   // alu.v(54)
    not (n184, n49) ;   // alu.v(54)
    not (n185, n48) ;   // alu.v(54)
    not (n186, n47) ;   // alu.v(54)
    not (n187, n46) ;   // alu.v(54)
    not (n188, n45) ;   // alu.v(54)
    not (n189, n44) ;   // alu.v(54)
    not (n190, n43) ;   // alu.v(54)
    not (n191, n42) ;   // alu.v(54)
    not (n192, n41) ;   // alu.v(54)
    not (n193, n40) ;   // alu.v(54)
    not (n194, n39) ;   // alu.v(54)
    not (n195, n38) ;   // alu.v(54)
    not (n196, n37) ;   // alu.v(54)
    not (n229, n100) ;   // alu.v(55)
    not (n230, n99) ;   // alu.v(55)
    not (n231, n98) ;   // alu.v(55)
    not (n232, n97) ;   // alu.v(55)
    not (n233, n96) ;   // alu.v(55)
    not (n234, n95) ;   // alu.v(55)
    not (n235, n94) ;   // alu.v(55)
    not (n236, n93) ;   // alu.v(55)
    not (n237, n92) ;   // alu.v(55)
    not (n238, n91) ;   // alu.v(55)
    not (n239, n90) ;   // alu.v(55)
    not (n240, n89) ;   // alu.v(55)
    not (n241, n88) ;   // alu.v(55)
    not (n242, n87) ;   // alu.v(55)
    not (n243, n86) ;   // alu.v(55)
    not (n244, n85) ;   // alu.v(55)
    not (n245, n84) ;   // alu.v(55)
    not (n246, n83) ;   // alu.v(55)
    not (n247, n82) ;   // alu.v(55)
    not (n248, n81) ;   // alu.v(55)
    not (n249, n80) ;   // alu.v(55)
    not (n250, n79) ;   // alu.v(55)
    not (n251, n78) ;   // alu.v(55)
    not (n252, n77) ;   // alu.v(55)
    not (n253, n76) ;   // alu.v(55)
    not (n254, n75) ;   // alu.v(55)
    not (n255, n74) ;   // alu.v(55)
    not (n256, n73) ;   // alu.v(55)
    not (n257, n72) ;   // alu.v(55)
    not (n258, n71) ;   // alu.v(55)
    not (n259, n70) ;   // alu.v(55)
    not (n260, n69) ;   // alu.v(55)
    not (n293, n132) ;   // alu.v(56)
    not (n294, n131) ;   // alu.v(56)
    not (n295, n130) ;   // alu.v(56)
    not (n296, n129) ;   // alu.v(56)
    not (n297, n128) ;   // alu.v(56)
    not (n298, n127) ;   // alu.v(56)
    not (n299, n126) ;   // alu.v(56)
    not (n300, n125) ;   // alu.v(56)
    not (n301, n124) ;   // alu.v(56)
    not (n302, n123) ;   // alu.v(56)
    not (n303, n122) ;   // alu.v(56)
    not (n304, n121) ;   // alu.v(56)
    not (n305, n120) ;   // alu.v(56)
    not (n306, n119) ;   // alu.v(56)
    not (n307, n118) ;   // alu.v(56)
    not (n308, n117) ;   // alu.v(56)
    not (n309, n116) ;   // alu.v(56)
    not (n310, n115) ;   // alu.v(56)
    not (n311, n114) ;   // alu.v(56)
    not (n312, n113) ;   // alu.v(56)
    not (n313, n112) ;   // alu.v(56)
    not (n314, n111) ;   // alu.v(56)
    not (n315, n110) ;   // alu.v(56)
    not (n316, n109) ;   // alu.v(56)
    not (n317, n108) ;   // alu.v(56)
    not (n318, n107) ;   // alu.v(56)
    not (n319, n106) ;   // alu.v(56)
    not (n320, n105) ;   // alu.v(56)
    not (n321, n104) ;   // alu.v(56)
    not (n322, n103) ;   // alu.v(56)
    not (n323, n102) ;   // alu.v(56)
    not (n324, n101) ;   // alu.v(56)
    not (n325, b[31]) ;   // alu.v(57)
    not (n326, b[30]) ;   // alu.v(57)
    not (n327, b[29]) ;   // alu.v(57)
    not (n328, b[28]) ;   // alu.v(57)
    not (n329, b[27]) ;   // alu.v(57)
    not (n330, b[26]) ;   // alu.v(57)
    not (n331, b[25]) ;   // alu.v(57)
    not (n332, b[24]) ;   // alu.v(57)
    not (n333, b[23]) ;   // alu.v(57)
    not (n334, b[22]) ;   // alu.v(57)
    not (n335, b[21]) ;   // alu.v(57)
    not (n336, b[20]) ;   // alu.v(57)
    not (n337, b[19]) ;   // alu.v(57)
    not (n338, b[18]) ;   // alu.v(57)
    not (n339, b[17]) ;   // alu.v(57)
    not (n340, b[16]) ;   // alu.v(57)
    not (n341, b[15]) ;   // alu.v(57)
    not (n342, b[14]) ;   // alu.v(57)
    not (n343, b[13]) ;   // alu.v(57)
    not (n344, b[12]) ;   // alu.v(57)
    not (n345, b[11]) ;   // alu.v(57)
    not (n346, b[10]) ;   // alu.v(57)
    not (n347, b[9]) ;   // alu.v(57)
    not (n348, b[8]) ;   // alu.v(57)
    not (n349, b[7]) ;   // alu.v(57)
    not (n350, b[6]) ;   // alu.v(57)
    not (n351, b[5]) ;   // alu.v(57)
    not (n352, b[4]) ;   // alu.v(57)
    not (n353, b[3]) ;   // alu.v(57)
    not (n354, b[2]) ;   // alu.v(57)
    not (n355, b[1]) ;   // alu.v(57)
    not (n356, b[0]) ;   // alu.v(57)
    Mux_3u_8u Mux_356 (.sel({op}), .data({n325, n293, n229, n165, 
            n132, n100, n68, n5}), .o(q[31]));   // alu.v(49)
    Mux_3u_8u Mux_357 (.sel({op}), .data({n326, n294, n230, n166, 
            n131, n99, n67, n6}), .o(q[30]));   // alu.v(49)
    Mux_3u_8u Mux_358 (.sel({op}), .data({n327, n295, n231, n167, 
            n130, n98, n66, n7}), .o(q[29]));   // alu.v(49)
    Mux_3u_8u Mux_359 (.sel({op}), .data({n328, n296, n232, n168, 
            n129, n97, n65, n8}), .o(q[28]));   // alu.v(49)
    Mux_3u_8u Mux_360 (.sel({op}), .data({n329, n297, n233, n169, 
            n128, n96, n64, n9}), .o(q[27]));   // alu.v(49)
    Mux_3u_8u Mux_361 (.sel({op}), .data({n330, n298, n234, n170, 
            n127, n95, n63, n10}), .o(q[26]));   // alu.v(49)
    Mux_3u_8u Mux_362 (.sel({op}), .data({n331, n299, n235, n171, 
            n126, n94, n62, n11}), .o(q[25]));   // alu.v(49)
    Mux_3u_8u Mux_363 (.sel({op}), .data({n332, n300, n236, n172, 
            n125, n93, n61, n12}), .o(q[24]));   // alu.v(49)
    Mux_3u_8u Mux_364 (.sel({op}), .data({n333, n301, n237, n173, 
            n124, n92, n60, n13}), .o(q[23]));   // alu.v(49)
    Mux_3u_8u Mux_365 (.sel({op}), .data({n334, n302, n238, n174, 
            n123, n91, n59, n14}), .o(q[22]));   // alu.v(49)
    Mux_3u_8u Mux_366 (.sel({op}), .data({n335, n303, n239, n175, 
            n122, n90, n58, n15}), .o(q[21]));   // alu.v(49)
    Mux_3u_8u Mux_367 (.sel({op}), .data({n336, n304, n240, n176, 
            n121, n89, n57, n16}), .o(q[20]));   // alu.v(49)
    Mux_3u_8u Mux_368 (.sel({op}), .data({n337, n305, n241, n177, 
            n120, n88, n56, n17}), .o(q[19]));   // alu.v(49)
    Mux_3u_8u Mux_369 (.sel({op}), .data({n338, n306, n242, n178, 
            n119, n87, n55, n18}), .o(q[18]));   // alu.v(49)
    Mux_3u_8u Mux_370 (.sel({op}), .data({n339, n307, n243, n179, 
            n118, n86, n54, n19}), .o(q[17]));   // alu.v(49)
    Mux_3u_8u Mux_371 (.sel({op}), .data({n340, n308, n244, n180, 
            n117, n85, n53, n20}), .o(q[16]));   // alu.v(49)
    Mux_3u_8u Mux_372 (.sel({op}), .data({n341, n309, n245, n181, 
            n116, n84, n52, n21}), .o(q[15]));   // alu.v(49)
    Mux_3u_8u Mux_373 (.sel({op}), .data({n342, n310, n246, n182, 
            n115, n83, n51, n22}), .o(q[14]));   // alu.v(49)
    Mux_3u_8u Mux_374 (.sel({op}), .data({n343, n311, n247, n183, 
            n114, n82, n50, n23}), .o(q[13]));   // alu.v(49)
    Mux_3u_8u Mux_375 (.sel({op}), .data({n344, n312, n248, n184, 
            n113, n81, n49, n24}), .o(q[12]));   // alu.v(49)
    Mux_3u_8u Mux_376 (.sel({op}), .data({n345, n313, n249, n185, 
            n112, n80, n48, n25}), .o(q[11]));   // alu.v(49)
    Mux_3u_8u Mux_377 (.sel({op}), .data({n346, n314, n250, n186, 
            n111, n79, n47, n26}), .o(q[10]));   // alu.v(49)
    Mux_3u_8u Mux_378 (.sel({op}), .data({n347, n315, n251, n187, 
            n110, n78, n46, n27}), .o(q[9]));   // alu.v(49)
    Mux_3u_8u Mux_379 (.sel({op}), .data({n348, n316, n252, n188, 
            n109, n77, n45, n28}), .o(q[8]));   // alu.v(49)
    Mux_3u_8u Mux_380 (.sel({op}), .data({n349, n317, n253, n189, 
            n108, n76, n44, n29}), .o(q[7]));   // alu.v(49)
    Mux_3u_8u Mux_381 (.sel({op}), .data({n350, n318, n254, n190, 
            n107, n75, n43, n30}), .o(q[6]));   // alu.v(49)
    Mux_3u_8u Mux_382 (.sel({op}), .data({n351, n319, n255, n191, 
            n106, n74, n42, n31}), .o(q[5]));   // alu.v(49)
    Mux_3u_8u Mux_383 (.sel({op}), .data({n352, n320, n256, n192, 
            n105, n73, n41, n32}), .o(q[4]));   // alu.v(49)
    Mux_3u_8u Mux_384 (.sel({op}), .data({n353, n321, n257, n193, 
            n104, n72, n40, n33}), .o(q[3]));   // alu.v(49)
    Mux_3u_8u Mux_385 (.sel({op}), .data({n354, n322, n258, n194, 
            n103, n71, n39, n34}), .o(q[2]));   // alu.v(49)
    Mux_3u_8u Mux_386 (.sel({op}), .data({n355, n323, n259, n195, 
            n102, n70, n38, n35}), .o(q[1]));   // alu.v(49)
    Mux_3u_8u Mux_387 (.sel({op}), .data({n356, n324, n260, n196, 
            n101, n69, n37, n36}), .o(q[0]));   // alu.v(49)
    
endmodule

//
// Verific Verilog Description of OPERATOR Select_6
//

module Select_6 (sel, data, o);
    input [5:0]sel;
    input [5:0]data;
    output o;
    assign o = |(sel & data);
    
endmodule

//
// Verific Verilog Description of PRIMITIVE VERIFIC_DLATCHRS
//

module VERIFIC_DLATCHRS (d, gate, s, r, q);
    input d;
    input gate;
    input s;
    input r;
    output q;
    reg q ;
    always @(gate or s or r or d) begin
        if (s) q = 1'b1;
        else if (r) q = 1'b0;
        else if (gate) q = d;
    end
    
endmodule

//
// Verific Verilog Description of module cond_calc
//

module cond_calc (cr, cc, n, z, c, v);   // execute.v(5)
    output cr;   // execute.v(9)
    input [3:0]cc;   // execute.v(6)
    input n;   // execute.v(7)
    input z;   // execute.v(7)
    input c;   // execute.v(7)
    input v;   // execute.v(7)
    
    
    wire n5, n7, n9, n11, n14, n17, n18, n19, n24, n27;
    
    not (n5, z) ;   // execute.v(14)
    not (n7, c) ;   // execute.v(16)
    not (n9, n) ;   // execute.v(18)
    not (n11, v) ;   // execute.v(20)
    and (n14, c, n5) ;   // execute.v(21)
    or (n17, n7, z) ;   // execute.v(22)
    xor (n18, n, v) ;   // execute.v(23)
    not (n19, n18) ;   // execute.v(23)
    and (n24, n5, n19) ;   // execute.v(25)
    or (n27, z, n18) ;   // execute.v(26)
    Mux_4u_16u Mux_27 (.sel({cc}), .data({2'b01, n27, n24, n18, n19, 
            n17, n14, n11, v, n9, n, n7, c, n5, z}), .o(cr));   // execute.v(12)
    
endmodule

//
// Verific Verilog Description of module status_register_adaptor
//

module status_register_adaptor (st, stwr, n, z, c, v, cc);   // execute.v(33)
    output [31:0]st;   // execute.v(37)
    output stwr;   // execute.v(38)
    input n;   // execute.v(34)
    input z;   // execute.v(34)
    input c;   // execute.v(34)
    input v;   // execute.v(34)
    input cc;   // execute.v(35)
    
    
    assign st[31] = 1'b0;   // execute.v(37)
    assign st[30] = 1'b0;   // execute.v(37)
    assign st[29] = 1'b0;   // execute.v(37)
    assign st[28] = 1'b0;   // execute.v(37)
    assign st[27] = 1'b0;   // execute.v(37)
    assign st[26] = 1'b0;   // execute.v(37)
    assign st[25] = 1'b0;   // execute.v(37)
    assign st[24] = 1'b0;   // execute.v(37)
    assign st[23] = 1'b0;   // execute.v(37)
    assign st[22] = 1'b0;   // execute.v(37)
    assign st[21] = 1'b0;   // execute.v(37)
    assign st[20] = 1'b0;   // execute.v(37)
    assign st[19] = 1'b0;   // execute.v(37)
    assign st[18] = 1'b0;   // execute.v(37)
    assign st[17] = 1'b0;   // execute.v(37)
    assign st[16] = 1'b0;   // execute.v(37)
    assign st[15] = 1'b0;   // execute.v(37)
    assign st[14] = 1'b0;   // execute.v(37)
    assign st[13] = 1'b0;   // execute.v(37)
    assign st[12] = 1'b0;   // execute.v(37)
    assign st[11] = 1'b0;   // execute.v(37)
    assign st[10] = 1'b0;   // execute.v(37)
    assign st[9] = 1'b0;   // execute.v(37)
    assign st[8] = 1'b0;   // execute.v(37)
    assign st[7] = 1'b0;   // execute.v(37)
    assign st[6] = 1'b0;   // execute.v(37)
    assign st[5] = 1'b0;   // execute.v(37)
    assign st[3] = n;   // execute.v(34)
    assign st[2] = z;   // execute.v(34)
    assign st[1] = c;   // execute.v(34)
    assign st[0] = v;   // execute.v(34)
    assign stwr = cc;   // execute.v(35)
    assign st[4] = 1'b0;
    
endmodule

//
// Verific Verilog Description of module execute_stage_passthrough
//

module execute_stage_passthrough (qm_a1, qm_a2, qm_r1_op, qm_r2_op, 
            qr_a1, qr_a2, qr_op, m_a1, m_a2, m_r1_op, m_r2_op, 
            r_a1, r_a2, r_op, clk, rst);   // execute.v(45)
    output [31:0]qm_a1;   // execute.v(54)
    output [31:0]qm_a2;   // execute.v(54)
    output [3:0]qm_r1_op;   // execute.v(55)
    output [3:0]qm_r2_op;   // execute.v(55)
    output [4:0]qr_a1;   // execute.v(57)
    output [4:0]qr_a2;   // execute.v(57)
    output [3:0]qr_op;   // execute.v(58)
    input [31:0]m_a1;   // execute.v(46)
    input [31:0]m_a2;   // execute.v(46)
    input [3:0]m_r1_op;   // execute.v(47)
    input [3:0]m_r2_op;   // execute.v(47)
    input [4:0]r_a1;   // execute.v(49)
    input [4:0]r_a2;   // execute.v(49)
    input [3:0]r_op;   // execute.v(50)
    input clk;   // execute.v(52)
    input rst;   // execute.v(52)
    
    
    VERIFIC_DFFRS i6 (.d(m_a1[30]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[30]));   // execute.v(67)
    VERIFIC_DFFRS i7 (.d(m_a1[29]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[29]));   // execute.v(67)
    VERIFIC_DFFRS i8 (.d(m_a1[28]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[28]));   // execute.v(67)
    VERIFIC_DFFRS i9 (.d(m_a1[27]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[27]));   // execute.v(67)
    VERIFIC_DFFRS i10 (.d(m_a1[26]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[26]));   // execute.v(67)
    VERIFIC_DFFRS i11 (.d(m_a1[25]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[25]));   // execute.v(67)
    VERIFIC_DFFRS i12 (.d(m_a1[24]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[24]));   // execute.v(67)
    VERIFIC_DFFRS i13 (.d(m_a1[23]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[23]));   // execute.v(67)
    VERIFIC_DFFRS i14 (.d(m_a1[22]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[22]));   // execute.v(67)
    VERIFIC_DFFRS i15 (.d(m_a1[21]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[21]));   // execute.v(67)
    VERIFIC_DFFRS i16 (.d(m_a1[20]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[20]));   // execute.v(67)
    VERIFIC_DFFRS i17 (.d(m_a1[19]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[19]));   // execute.v(67)
    VERIFIC_DFFRS i18 (.d(m_a1[18]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[18]));   // execute.v(67)
    VERIFIC_DFFRS i19 (.d(m_a1[17]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[17]));   // execute.v(67)
    VERIFIC_DFFRS i20 (.d(m_a1[16]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[16]));   // execute.v(67)
    VERIFIC_DFFRS i21 (.d(m_a1[15]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[15]));   // execute.v(67)
    VERIFIC_DFFRS i22 (.d(m_a1[14]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[14]));   // execute.v(67)
    VERIFIC_DFFRS i23 (.d(m_a1[13]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[13]));   // execute.v(67)
    VERIFIC_DFFRS i24 (.d(m_a1[12]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[12]));   // execute.v(67)
    VERIFIC_DFFRS i25 (.d(m_a1[11]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[11]));   // execute.v(67)
    VERIFIC_DFFRS i26 (.d(m_a1[10]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[10]));   // execute.v(67)
    VERIFIC_DFFRS i27 (.d(m_a1[9]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[9]));   // execute.v(67)
    VERIFIC_DFFRS i28 (.d(m_a1[8]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[8]));   // execute.v(67)
    VERIFIC_DFFRS i29 (.d(m_a1[7]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[7]));   // execute.v(67)
    VERIFIC_DFFRS i30 (.d(m_a1[6]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[6]));   // execute.v(67)
    VERIFIC_DFFRS i31 (.d(m_a1[5]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[5]));   // execute.v(67)
    VERIFIC_DFFRS i32 (.d(m_a1[4]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[4]));   // execute.v(67)
    VERIFIC_DFFRS i33 (.d(m_a1[3]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[3]));   // execute.v(67)
    VERIFIC_DFFRS i34 (.d(m_a1[2]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[2]));   // execute.v(67)
    VERIFIC_DFFRS i35 (.d(m_a1[1]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[1]));   // execute.v(67)
    VERIFIC_DFFRS i36 (.d(m_a1[0]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[0]));   // execute.v(67)
    VERIFIC_DFFRS i37 (.d(m_a2[31]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[31]));   // execute.v(67)
    VERIFIC_DFFRS i38 (.d(m_a2[30]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[30]));   // execute.v(67)
    VERIFIC_DFFRS i39 (.d(m_a2[29]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[29]));   // execute.v(67)
    VERIFIC_DFFRS i40 (.d(m_a2[28]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[28]));   // execute.v(67)
    VERIFIC_DFFRS i41 (.d(m_a2[27]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[27]));   // execute.v(67)
    VERIFIC_DFFRS i42 (.d(m_a2[26]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[26]));   // execute.v(67)
    VERIFIC_DFFRS i43 (.d(m_a2[25]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[25]));   // execute.v(67)
    VERIFIC_DFFRS i44 (.d(m_a2[24]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[24]));   // execute.v(67)
    VERIFIC_DFFRS i45 (.d(m_a2[23]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[23]));   // execute.v(67)
    VERIFIC_DFFRS i46 (.d(m_a2[22]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[22]));   // execute.v(67)
    VERIFIC_DFFRS i47 (.d(m_a2[21]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[21]));   // execute.v(67)
    VERIFIC_DFFRS i48 (.d(m_a2[20]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[20]));   // execute.v(67)
    VERIFIC_DFFRS i49 (.d(m_a2[19]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[19]));   // execute.v(67)
    VERIFIC_DFFRS i50 (.d(m_a2[18]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[18]));   // execute.v(67)
    VERIFIC_DFFRS i51 (.d(m_a2[17]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[17]));   // execute.v(67)
    VERIFIC_DFFRS i52 (.d(m_a2[16]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[16]));   // execute.v(67)
    VERIFIC_DFFRS i53 (.d(m_a2[15]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[15]));   // execute.v(67)
    VERIFIC_DFFRS i54 (.d(m_a2[14]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[14]));   // execute.v(67)
    VERIFIC_DFFRS i55 (.d(m_a2[13]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[13]));   // execute.v(67)
    VERIFIC_DFFRS i56 (.d(m_a2[12]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[12]));   // execute.v(67)
    VERIFIC_DFFRS i57 (.d(m_a2[11]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[11]));   // execute.v(67)
    VERIFIC_DFFRS i58 (.d(m_a2[10]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[10]));   // execute.v(67)
    VERIFIC_DFFRS i59 (.d(m_a2[9]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[9]));   // execute.v(67)
    VERIFIC_DFFRS i60 (.d(m_a2[8]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[8]));   // execute.v(67)
    VERIFIC_DFFRS i61 (.d(m_a2[7]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[7]));   // execute.v(67)
    VERIFIC_DFFRS i62 (.d(m_a2[6]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[6]));   // execute.v(67)
    VERIFIC_DFFRS i63 (.d(m_a2[5]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[5]));   // execute.v(67)
    VERIFIC_DFFRS i64 (.d(m_a2[4]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[4]));   // execute.v(67)
    VERIFIC_DFFRS i65 (.d(m_a2[3]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[3]));   // execute.v(67)
    VERIFIC_DFFRS i66 (.d(m_a2[2]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[2]));   // execute.v(67)
    VERIFIC_DFFRS i67 (.d(m_a2[1]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[1]));   // execute.v(67)
    VERIFIC_DFFRS i68 (.d(m_a2[0]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a2[0]));   // execute.v(67)
    VERIFIC_DFFRS i69 (.d(m_r1_op[3]), .clk(clk), .s(1'b0), .r(rst), 
            .q(qm_r1_op[3]));   // execute.v(67)
    VERIFIC_DFFRS i70 (.d(m_r1_op[2]), .clk(clk), .s(1'b0), .r(rst), 
            .q(qm_r1_op[2]));   // execute.v(67)
    VERIFIC_DFFRS i71 (.d(m_r1_op[1]), .clk(clk), .s(1'b0), .r(rst), 
            .q(qm_r1_op[1]));   // execute.v(67)
    VERIFIC_DFFRS i72 (.d(m_r1_op[0]), .clk(clk), .s(1'b0), .r(rst), 
            .q(qm_r1_op[0]));   // execute.v(67)
    VERIFIC_DFFRS i73 (.d(m_r2_op[3]), .clk(clk), .s(1'b0), .r(rst), 
            .q(qm_r2_op[3]));   // execute.v(67)
    VERIFIC_DFFRS i74 (.d(m_r2_op[2]), .clk(clk), .s(1'b0), .r(rst), 
            .q(qm_r2_op[2]));   // execute.v(67)
    VERIFIC_DFFRS i75 (.d(m_r2_op[1]), .clk(clk), .s(1'b0), .r(rst), 
            .q(qm_r2_op[1]));   // execute.v(67)
    VERIFIC_DFFRS i76 (.d(m_r2_op[0]), .clk(clk), .s(1'b0), .r(rst), 
            .q(qm_r2_op[0]));   // execute.v(67)
    VERIFIC_DFFRS i77 (.d(r_a1[4]), .clk(clk), .s(1'b0), .r(rst), .q(qr_a1[4]));   // execute.v(67)
    VERIFIC_DFFRS i78 (.d(r_a1[3]), .clk(clk), .s(1'b0), .r(rst), .q(qr_a1[3]));   // execute.v(67)
    VERIFIC_DFFRS i79 (.d(r_a1[2]), .clk(clk), .s(1'b0), .r(rst), .q(qr_a1[2]));   // execute.v(67)
    VERIFIC_DFFRS i80 (.d(r_a1[1]), .clk(clk), .s(1'b0), .r(rst), .q(qr_a1[1]));   // execute.v(67)
    VERIFIC_DFFRS i81 (.d(r_a1[0]), .clk(clk), .s(1'b0), .r(rst), .q(qr_a1[0]));   // execute.v(67)
    VERIFIC_DFFRS i82 (.d(r_a2[4]), .clk(clk), .s(1'b0), .r(rst), .q(qr_a2[4]));   // execute.v(67)
    VERIFIC_DFFRS i83 (.d(r_a2[3]), .clk(clk), .s(1'b0), .r(rst), .q(qr_a2[3]));   // execute.v(67)
    VERIFIC_DFFRS i84 (.d(r_a2[2]), .clk(clk), .s(1'b0), .r(rst), .q(qr_a2[2]));   // execute.v(67)
    VERIFIC_DFFRS i85 (.d(r_a2[1]), .clk(clk), .s(1'b0), .r(rst), .q(qr_a2[1]));   // execute.v(67)
    VERIFIC_DFFRS i86 (.d(r_a2[0]), .clk(clk), .s(1'b0), .r(rst), .q(qr_a2[0]));   // execute.v(67)
    VERIFIC_DFFRS i87 (.d(r_op[3]), .clk(clk), .s(1'b0), .r(rst), .q(qr_op[3]));   // execute.v(67)
    VERIFIC_DFFRS i88 (.d(r_op[2]), .clk(clk), .s(1'b0), .r(rst), .q(qr_op[2]));   // execute.v(67)
    VERIFIC_DFFRS i89 (.d(r_op[1]), .clk(clk), .s(1'b0), .r(rst), .q(qr_op[1]));   // execute.v(67)
    VERIFIC_DFFRS i90 (.d(r_op[0]), .clk(clk), .s(1'b0), .r(rst), .q(qr_op[0]));   // execute.v(67)
    VERIFIC_DFFRS i5 (.d(m_a1[31]), .clk(clk), .s(1'b0), .r(rst), .q(qm_a1[31]));   // execute.v(67)
    
endmodule

//
// Verific Verilog Description of module memory_op
//

module memory_op (m1, m2, ram_w_addr, ram_r_addr, ram_w, ram_r, 
            ram_w_line, sys_w_addr, sys_r_addr, sys_w, sys_r, sys_w_line, 
            r1, r2, a1, a2, r1_op, r2_op, ram_r_line, sys_r_line, 
            proceed, clk, rst);   // memory_op.v(28)
    output [31:0]m1;   // memory_op.v(40)
    output [31:0]m2;   // memory_op.v(40)
    output [31:0]ram_w_addr;   // memory_op.v(42)
    output [31:0]ram_r_addr;   // memory_op.v(43)
    output ram_w;   // memory_op.v(47)
    output ram_r;   // memory_op.v(47)
    output [31:0]ram_w_line;   // memory_op.v(45)
    output [31:0]sys_w_addr;   // memory_op.v(42)
    output [31:0]sys_r_addr;   // memory_op.v(43)
    output sys_w;   // memory_op.v(47)
    output sys_r;   // memory_op.v(47)
    output [31:0]sys_w_line;   // memory_op.v(45)
    input [31:0]r1;   // memory_op.v(29)
    input [31:0]r2;   // memory_op.v(29)
    input [31:0]a1;   // memory_op.v(30)
    input [31:0]a2;   // memory_op.v(30)
    input [3:0]r1_op;   // memory_op.v(32)
    input [3:0]r2_op;   // memory_op.v(32)
    input [31:0]ram_r_line;   // memory_op.v(34)
    input [31:0]sys_r_line;   // memory_op.v(34)
    input proceed;   // memory_op.v(36)
    input clk;   // memory_op.v(38)
    input rst;   // memory_op.v(38)
    
    wire [3:0]r1_op_inner;   // memory_op.v(49)
    wire [3:0]r2_op_inner;   // memory_op.v(49)
    wire [31:0]r1_inner;   // memory_op.v(54)
    wire [31:0]r2_inner;   // memory_op.v(54)
    wire [2:0]m1_select;   // memory_op.v(56)
    wire [2:0]m2_select;   // memory_op.v(56)
    
    wire n12, n13, n14, n15, n16, n19, n20, n21, n22, n23, 
        n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, 
        n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
        n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, 
        n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
        n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, 
        n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, 
        n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, 
        n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, 
        n104, n105, n106, n107, n108, n109, n110, n111, n112, 
        n113, n114, n115, n116, n117, n118, n119, n120, n121, 
        n122, n123, n124, n125, n126, n127, n128, n129, n130, 
        n131, n132, n133, n134, n135, n136, n137, n138, n139, 
        n140, n141, n142, n143, n144, n145, n146, n147, n148, 
        n149, n182, n183, n184, n185, n186, n189, n190, n191, 
        n192, n193, n194, n195, n196, n197, n198, n199, n200, 
        n201, n202, n203, n204, n205, n206, n207, n208, n209, 
        n210, n211, n212, n213, n214, n215, n216, n217, n218, 
        n219, n220, n221, n222, n223, n224, n225, n226, n227, 
        n228, n229, n230, n231, n232, n233, n234, n235, n236, 
        n237, n238, n239, n240, n241, n242, n243, n244, n245, 
        n246, n247, n248, n249, n250, n251, n252, n253, n254, 
        n255, n256, n257, n258, n259, n260, n261, n262, n263, 
        n264, n265, n266, n267, n268, n269, n270, n271, n272, 
        n273, n274, n275, n276, n277, n278, n279, n280, n281, 
        n282, n283, n284, n285, n286, n287, n288, n289, n290, 
        n291, n292, n293, n294, n295, n296, n297, n298, n299, 
        n300, n301, n302, n303, n304, n305, n306, n307, n308, 
        n309, n310, n311, n312, n313, n314, n315, n316, n317, 
        n318, n319, n353, n354, n355, n356, n357, n358, n359, 
        n360, n361, n362, n363, n364, n365, n366, n367, n368, 
        n369, n370, n371, n372, n373, n374, n375, n376, n377, 
        n378, n379, n380, n381, n382, n383, n384, n385, n386, 
        n387, n388, n389, n390, n391, n392, n393, n394, n395, 
        n396, n397, n398, n399, n400, n401, n402, n403, n404, 
        n405, n406, n407, n408, n409, n410, n411, n412, n413, 
        n414, n415, n416, n417, n418, n419, n420, n421, n422, 
        n423, n424, n425, n426, n427, n428, n429, n430, n431, 
        n432, n433, n434, n435, n436, n437, n438, n439, n440, 
        n441, n442, n443, n444, n445, n446, n447, n448, n449, 
        n450, n451, n452, n453, n454, n455, n456, n457, n458, 
        n459, n460, n461, n462, n463, n464, n465, n466, n467, 
        n468, n469, n470, n471, n472, n473, n474, n475, n476, 
        n477, n478, n479, n480, n481, n482, n483, n484, n485, 
        n486, n487, n488, n489, n490, n491, n492, n493, n494, 
        n495, n496, n497, n498, n499, n500, n501, n502, n503, 
        n504, n505, n506, n507, n508, n509, n510, n511, n512, 
        n513, n514, n515, n516, n517, n518, n519, n520, n521, 
        n522, n523, n524, n525, n526, n527, n528, n529, n530, 
        n531, n532, n533, n534, n535, n536, n537, n538, n539, 
        n540, n541, n542, n543, n544, n545, n546, n547, n548, 
        n549, n550, n551, n552, n553, n554, n555, n556, n557, 
        n558, n559, n560, n561, n562, n563, n564, n565, n566, 
        n567, n568, n569, n570, n571, n572, n573, n574, n575, 
        n576, n577, n578, n579, n580, n581, n582, n583, n584, 
        n585, n586, n587, n588, n589, n590, n591, n592, n593, 
        n594, n595, n596, n597, n598, n599, n600, n601, n602, 
        n603, n604, n605, n606, n607, n608, n609, n610, n611, 
        n612, n613, n614, n615, n616, n617, n618, n619, n620, 
        n621, n622, n623, n624, n625, n626, n627, n628, n629, 
        n630, n631, n632, n633, n634, n635, n636, n637, n638, 
        n639, n640, n641, n642, n643, n644, n645, n646, n647, 
        n648, n649, n650, n651, n652, n653, n654, n655, n656, 
        n657, n658, n659, n660, n661, n662, n663, n664, n665, 
        n666, n667, n668, n669, n670, n671, n672, n673, n674, 
        n675, n676, n677, n678, n679, n680, n681, n682, n683, 
        n684, n685, n686, n687, n688, n689, n690, n691, n692, 
        n693, n694, n695, n696, n697, n698, n699, n700, n701, 
        n702, n703, n704, n705, n706, n707, n708, n709, n710, 
        n711, n712, n713, n714, n715, n716, n717, n718, n719, 
        n720, n721, n722, n723, n724, n725, n726, n727, n728, 
        n729, n730, n731, n732, n733, n734, n735, n736, n737, 
        n738, n739, n740, n741, n742, n743, n744, n745, n746, 
        n747, n748, n749, n750;
    
    assign r1_op_inner[3] = proceed ? r1_op[3] : 1'b0;   // memory_op.v(51)
    assign r1_op_inner[2] = proceed ? r1_op[2] : 1'b0;   // memory_op.v(51)
    assign r1_op_inner[1] = proceed ? r1_op[1] : 1'b0;   // memory_op.v(51)
    assign r1_op_inner[0] = proceed ? r1_op[0] : 1'b0;   // memory_op.v(51)
    assign r2_op_inner[3] = proceed ? r2_op[3] : 1'b0;   // memory_op.v(52)
    assign r2_op_inner[2] = proceed ? r2_op[2] : 1'b0;   // memory_op.v(52)
    assign r2_op_inner[1] = proceed ? r2_op[1] : 1'b0;   // memory_op.v(52)
    assign r2_op_inner[0] = proceed ? r2_op[0] : 1'b0;   // memory_op.v(52)
    nor (n12, m1_select[2], m1_select[1], m1_select[0]) ;   // memory_op.v(57)
    not (n13, m1_select[0]) ;   // memory_op.v(57)
    nor (n14, m1_select[2], m1_select[1], n13) ;   // memory_op.v(57)
    not (n15, m1_select[1]) ;   // memory_op.v(57)
    nor (n16, m1_select[2], n15, m1_select[0]) ;   // memory_op.v(57)
    nor (n19, m1_select[2], n15, n13) ;   // memory_op.v(57)
    not (n20, m1_select[2]) ;   // memory_op.v(57)
    nor (n21, n20, m1_select[1], m1_select[0]) ;   // memory_op.v(57)
    assign n22 = n21 ? sys_r_line[31] : 1'b1;   // memory_op.v(57)
    assign n23 = n21 ? sys_r_line[30] : 1'b0;   // memory_op.v(57)
    assign n24 = n21 ? sys_r_line[29] : 1'b1;   // memory_op.v(57)
    assign n25 = n21 ? sys_r_line[28] : 1'b0;   // memory_op.v(57)
    assign n26 = n21 ? sys_r_line[27] : 1'b1;   // memory_op.v(57)
    assign n27 = n21 ? sys_r_line[26] : 1'b0;   // memory_op.v(57)
    assign n28 = n21 ? sys_r_line[25] : 1'b1;   // memory_op.v(57)
    assign n29 = n21 ? sys_r_line[24] : 1'b0;   // memory_op.v(57)
    assign n30 = n21 ? sys_r_line[23] : 1'b1;   // memory_op.v(57)
    assign n31 = n21 ? sys_r_line[22] : 1'b0;   // memory_op.v(57)
    assign n32 = n21 ? sys_r_line[21] : 1'b1;   // memory_op.v(57)
    assign n33 = n21 ? sys_r_line[20] : 1'b0;   // memory_op.v(57)
    assign n34 = n21 ? sys_r_line[19] : 1'b1;   // memory_op.v(57)
    assign n35 = n21 ? sys_r_line[18] : 1'b0;   // memory_op.v(57)
    assign n36 = n21 ? sys_r_line[17] : 1'b1;   // memory_op.v(57)
    assign n37 = n21 ? sys_r_line[16] : 1'b0;   // memory_op.v(57)
    assign n38 = n21 ? sys_r_line[15] : 1'b1;   // memory_op.v(57)
    assign n39 = n21 ? sys_r_line[14] : 1'b0;   // memory_op.v(57)
    assign n40 = n21 ? sys_r_line[13] : 1'b1;   // memory_op.v(57)
    assign n41 = n21 ? sys_r_line[12] : 1'b0;   // memory_op.v(57)
    assign n42 = n21 ? sys_r_line[11] : 1'b1;   // memory_op.v(57)
    assign n43 = n21 ? sys_r_line[10] : 1'b0;   // memory_op.v(57)
    assign n44 = n21 ? sys_r_line[9] : 1'b1;   // memory_op.v(57)
    assign n45 = n21 ? sys_r_line[8] : 1'b0;   // memory_op.v(57)
    assign n46 = n21 ? sys_r_line[7] : 1'b1;   // memory_op.v(57)
    assign n47 = n21 ? sys_r_line[6] : 1'b0;   // memory_op.v(57)
    assign n48 = n21 ? sys_r_line[5] : 1'b1;   // memory_op.v(57)
    assign n49 = n21 ? sys_r_line[4] : 1'b0;   // memory_op.v(57)
    assign n50 = n21 ? sys_r_line[3] : 1'b1;   // memory_op.v(57)
    assign n51 = n21 ? sys_r_line[2] : 1'b0;   // memory_op.v(57)
    assign n52 = n21 ? sys_r_line[1] : 1'b1;   // memory_op.v(57)
    assign n53 = n21 ? sys_r_line[0] : 1'b0;   // memory_op.v(57)
    assign n54 = n19 ? ram_r_line[31] : n22;   // memory_op.v(57)
    assign n55 = n19 ? ram_r_line[30] : n23;   // memory_op.v(57)
    assign n56 = n19 ? ram_r_line[29] : n24;   // memory_op.v(57)
    assign n57 = n19 ? ram_r_line[28] : n25;   // memory_op.v(57)
    assign n58 = n19 ? ram_r_line[27] : n26;   // memory_op.v(57)
    assign n59 = n19 ? ram_r_line[26] : n27;   // memory_op.v(57)
    assign n60 = n19 ? ram_r_line[25] : n28;   // memory_op.v(57)
    assign n61 = n19 ? ram_r_line[24] : n29;   // memory_op.v(57)
    assign n62 = n19 ? ram_r_line[23] : n30;   // memory_op.v(57)
    assign n63 = n19 ? ram_r_line[22] : n31;   // memory_op.v(57)
    assign n64 = n19 ? ram_r_line[21] : n32;   // memory_op.v(57)
    assign n65 = n19 ? ram_r_line[20] : n33;   // memory_op.v(57)
    assign n66 = n19 ? ram_r_line[19] : n34;   // memory_op.v(57)
    assign n67 = n19 ? ram_r_line[18] : n35;   // memory_op.v(57)
    assign n68 = n19 ? ram_r_line[17] : n36;   // memory_op.v(57)
    assign n69 = n19 ? ram_r_line[16] : n37;   // memory_op.v(57)
    assign n70 = n19 ? ram_r_line[15] : n38;   // memory_op.v(57)
    assign n71 = n19 ? ram_r_line[14] : n39;   // memory_op.v(57)
    assign n72 = n19 ? ram_r_line[13] : n40;   // memory_op.v(57)
    assign n73 = n19 ? ram_r_line[12] : n41;   // memory_op.v(57)
    assign n74 = n19 ? ram_r_line[11] : n42;   // memory_op.v(57)
    assign n75 = n19 ? ram_r_line[10] : n43;   // memory_op.v(57)
    assign n76 = n19 ? ram_r_line[9] : n44;   // memory_op.v(57)
    assign n77 = n19 ? ram_r_line[8] : n45;   // memory_op.v(57)
    assign n78 = n19 ? ram_r_line[7] : n46;   // memory_op.v(57)
    assign n79 = n19 ? ram_r_line[6] : n47;   // memory_op.v(57)
    assign n80 = n19 ? ram_r_line[5] : n48;   // memory_op.v(57)
    assign n81 = n19 ? ram_r_line[4] : n49;   // memory_op.v(57)
    assign n82 = n19 ? ram_r_line[3] : n50;   // memory_op.v(57)
    assign n83 = n19 ? ram_r_line[2] : n51;   // memory_op.v(57)
    assign n84 = n19 ? ram_r_line[1] : n52;   // memory_op.v(57)
    assign n85 = n19 ? ram_r_line[0] : n53;   // memory_op.v(57)
    assign n86 = n16 ? r2_inner[31] : n54;   // memory_op.v(57)
    assign n87 = n16 ? r2_inner[30] : n55;   // memory_op.v(57)
    assign n88 = n16 ? r2_inner[29] : n56;   // memory_op.v(57)
    assign n89 = n16 ? r2_inner[28] : n57;   // memory_op.v(57)
    assign n90 = n16 ? r2_inner[27] : n58;   // memory_op.v(57)
    assign n91 = n16 ? r2_inner[26] : n59;   // memory_op.v(57)
    assign n92 = n16 ? r2_inner[25] : n60;   // memory_op.v(57)
    assign n93 = n16 ? r2_inner[24] : n61;   // memory_op.v(57)
    assign n94 = n16 ? r2_inner[23] : n62;   // memory_op.v(57)
    assign n95 = n16 ? r2_inner[22] : n63;   // memory_op.v(57)
    assign n96 = n16 ? r2_inner[21] : n64;   // memory_op.v(57)
    assign n97 = n16 ? r2_inner[20] : n65;   // memory_op.v(57)
    assign n98 = n16 ? r2_inner[19] : n66;   // memory_op.v(57)
    assign n99 = n16 ? r2_inner[18] : n67;   // memory_op.v(57)
    assign n100 = n16 ? r2_inner[17] : n68;   // memory_op.v(57)
    assign n101 = n16 ? r2_inner[16] : n69;   // memory_op.v(57)
    assign n102 = n16 ? r2_inner[15] : n70;   // memory_op.v(57)
    assign n103 = n16 ? r2_inner[14] : n71;   // memory_op.v(57)
    assign n104 = n16 ? r2_inner[13] : n72;   // memory_op.v(57)
    assign n105 = n16 ? r2_inner[12] : n73;   // memory_op.v(57)
    assign n106 = n16 ? r2_inner[11] : n74;   // memory_op.v(57)
    assign n107 = n16 ? r2_inner[10] : n75;   // memory_op.v(57)
    assign n108 = n16 ? r2_inner[9] : n76;   // memory_op.v(57)
    assign n109 = n16 ? r2_inner[8] : n77;   // memory_op.v(57)
    assign n110 = n16 ? r2_inner[7] : n78;   // memory_op.v(57)
    assign n111 = n16 ? r2_inner[6] : n79;   // memory_op.v(57)
    assign n112 = n16 ? r2_inner[5] : n80;   // memory_op.v(57)
    assign n113 = n16 ? r2_inner[4] : n81;   // memory_op.v(57)
    assign n114 = n16 ? r2_inner[3] : n82;   // memory_op.v(57)
    assign n115 = n16 ? r2_inner[2] : n83;   // memory_op.v(57)
    assign n116 = n16 ? r2_inner[1] : n84;   // memory_op.v(57)
    assign n117 = n16 ? r2_inner[0] : n85;   // memory_op.v(57)
    assign n118 = n14 ? r1_inner[31] : n86;   // memory_op.v(57)
    assign n119 = n14 ? r1_inner[30] : n87;   // memory_op.v(57)
    assign n120 = n14 ? r1_inner[29] : n88;   // memory_op.v(57)
    assign n121 = n14 ? r1_inner[28] : n89;   // memory_op.v(57)
    assign n122 = n14 ? r1_inner[27] : n90;   // memory_op.v(57)
    assign n123 = n14 ? r1_inner[26] : n91;   // memory_op.v(57)
    assign n124 = n14 ? r1_inner[25] : n92;   // memory_op.v(57)
    assign n125 = n14 ? r1_inner[24] : n93;   // memory_op.v(57)
    assign n126 = n14 ? r1_inner[23] : n94;   // memory_op.v(57)
    assign n127 = n14 ? r1_inner[22] : n95;   // memory_op.v(57)
    assign n128 = n14 ? r1_inner[21] : n96;   // memory_op.v(57)
    assign n129 = n14 ? r1_inner[20] : n97;   // memory_op.v(57)
    assign n130 = n14 ? r1_inner[19] : n98;   // memory_op.v(57)
    assign n131 = n14 ? r1_inner[18] : n99;   // memory_op.v(57)
    assign n132 = n14 ? r1_inner[17] : n100;   // memory_op.v(57)
    assign n133 = n14 ? r1_inner[16] : n101;   // memory_op.v(57)
    assign n134 = n14 ? r1_inner[15] : n102;   // memory_op.v(57)
    assign n135 = n14 ? r1_inner[14] : n103;   // memory_op.v(57)
    assign n136 = n14 ? r1_inner[13] : n104;   // memory_op.v(57)
    assign n137 = n14 ? r1_inner[12] : n105;   // memory_op.v(57)
    assign n138 = n14 ? r1_inner[11] : n106;   // memory_op.v(57)
    assign n139 = n14 ? r1_inner[10] : n107;   // memory_op.v(57)
    assign n140 = n14 ? r1_inner[9] : n108;   // memory_op.v(57)
    assign n141 = n14 ? r1_inner[8] : n109;   // memory_op.v(57)
    assign n142 = n14 ? r1_inner[7] : n110;   // memory_op.v(57)
    assign n143 = n14 ? r1_inner[6] : n111;   // memory_op.v(57)
    assign n144 = n14 ? r1_inner[5] : n112;   // memory_op.v(57)
    assign n145 = n14 ? r1_inner[4] : n113;   // memory_op.v(57)
    assign n146 = n14 ? r1_inner[3] : n114;   // memory_op.v(57)
    assign n147 = n14 ? r1_inner[2] : n115;   // memory_op.v(57)
    assign n148 = n14 ? r1_inner[1] : n116;   // memory_op.v(57)
    assign n149 = n14 ? r1_inner[0] : n117;   // memory_op.v(57)
    assign m1[31] = n12 ? 1'b0 : n118;   // memory_op.v(57)
    assign m1[30] = n12 ? 1'b0 : n119;   // memory_op.v(57)
    assign m1[29] = n12 ? 1'b0 : n120;   // memory_op.v(57)
    assign m1[28] = n12 ? 1'b0 : n121;   // memory_op.v(57)
    assign m1[27] = n12 ? 1'b0 : n122;   // memory_op.v(57)
    assign m1[26] = n12 ? 1'b0 : n123;   // memory_op.v(57)
    assign m1[25] = n12 ? 1'b0 : n124;   // memory_op.v(57)
    assign m1[24] = n12 ? 1'b0 : n125;   // memory_op.v(57)
    assign m1[23] = n12 ? 1'b0 : n126;   // memory_op.v(57)
    assign m1[22] = n12 ? 1'b0 : n127;   // memory_op.v(57)
    assign m1[21] = n12 ? 1'b0 : n128;   // memory_op.v(57)
    assign m1[20] = n12 ? 1'b0 : n129;   // memory_op.v(57)
    assign m1[19] = n12 ? 1'b0 : n130;   // memory_op.v(57)
    assign m1[18] = n12 ? 1'b0 : n131;   // memory_op.v(57)
    assign m1[17] = n12 ? 1'b0 : n132;   // memory_op.v(57)
    assign m1[16] = n12 ? 1'b0 : n133;   // memory_op.v(57)
    assign m1[15] = n12 ? 1'b0 : n134;   // memory_op.v(57)
    assign m1[14] = n12 ? 1'b0 : n135;   // memory_op.v(57)
    assign m1[13] = n12 ? 1'b0 : n136;   // memory_op.v(57)
    assign m1[12] = n12 ? 1'b0 : n137;   // memory_op.v(57)
    assign m1[11] = n12 ? 1'b0 : n138;   // memory_op.v(57)
    assign m1[10] = n12 ? 1'b0 : n139;   // memory_op.v(57)
    assign m1[9] = n12 ? 1'b0 : n140;   // memory_op.v(57)
    assign m1[8] = n12 ? 1'b0 : n141;   // memory_op.v(57)
    assign m1[7] = n12 ? 1'b0 : n142;   // memory_op.v(57)
    assign m1[6] = n12 ? 1'b0 : n143;   // memory_op.v(57)
    assign m1[5] = n12 ? 1'b0 : n144;   // memory_op.v(57)
    assign m1[4] = n12 ? 1'b0 : n145;   // memory_op.v(57)
    assign m1[3] = n12 ? 1'b0 : n146;   // memory_op.v(57)
    assign m1[2] = n12 ? 1'b0 : n147;   // memory_op.v(57)
    assign m1[1] = n12 ? 1'b0 : n148;   // memory_op.v(57)
    assign m1[0] = n12 ? 1'b0 : n149;   // memory_op.v(57)
    nor (n182, m2_select[2], m2_select[1], m2_select[0]) ;   // memory_op.v(58)
    not (n183, m2_select[0]) ;   // memory_op.v(58)
    nor (n184, m2_select[2], m2_select[1], n183) ;   // memory_op.v(58)
    not (n185, m2_select[1]) ;   // memory_op.v(58)
    nor (n186, m2_select[2], n185, m2_select[0]) ;   // memory_op.v(58)
    nor (n189, m2_select[2], n185, n183) ;   // memory_op.v(58)
    not (n190, m2_select[2]) ;   // memory_op.v(58)
    nor (n191, n190, m2_select[1], m2_select[0]) ;   // memory_op.v(58)
    assign n192 = n191 ? sys_r_line[31] : 1'b1;   // memory_op.v(58)
    assign n193 = n191 ? sys_r_line[30] : 1'b0;   // memory_op.v(58)
    assign n194 = n191 ? sys_r_line[29] : 1'b1;   // memory_op.v(58)
    assign n195 = n191 ? sys_r_line[28] : 1'b0;   // memory_op.v(58)
    assign n196 = n191 ? sys_r_line[27] : 1'b1;   // memory_op.v(58)
    assign n197 = n191 ? sys_r_line[26] : 1'b0;   // memory_op.v(58)
    assign n198 = n191 ? sys_r_line[25] : 1'b1;   // memory_op.v(58)
    assign n199 = n191 ? sys_r_line[24] : 1'b0;   // memory_op.v(58)
    assign n200 = n191 ? sys_r_line[23] : 1'b1;   // memory_op.v(58)
    assign n201 = n191 ? sys_r_line[22] : 1'b0;   // memory_op.v(58)
    assign n202 = n191 ? sys_r_line[21] : 1'b1;   // memory_op.v(58)
    assign n203 = n191 ? sys_r_line[20] : 1'b0;   // memory_op.v(58)
    assign n204 = n191 ? sys_r_line[19] : 1'b1;   // memory_op.v(58)
    assign n205 = n191 ? sys_r_line[18] : 1'b0;   // memory_op.v(58)
    assign n206 = n191 ? sys_r_line[17] : 1'b1;   // memory_op.v(58)
    assign n207 = n191 ? sys_r_line[16] : 1'b0;   // memory_op.v(58)
    assign n208 = n191 ? sys_r_line[15] : 1'b1;   // memory_op.v(58)
    assign n209 = n191 ? sys_r_line[14] : 1'b0;   // memory_op.v(58)
    assign n210 = n191 ? sys_r_line[13] : 1'b1;   // memory_op.v(58)
    assign n211 = n191 ? sys_r_line[12] : 1'b0;   // memory_op.v(58)
    assign n212 = n191 ? sys_r_line[11] : 1'b1;   // memory_op.v(58)
    assign n213 = n191 ? sys_r_line[10] : 1'b0;   // memory_op.v(58)
    assign n214 = n191 ? sys_r_line[9] : 1'b1;   // memory_op.v(58)
    assign n215 = n191 ? sys_r_line[8] : 1'b0;   // memory_op.v(58)
    assign n216 = n191 ? sys_r_line[7] : 1'b1;   // memory_op.v(58)
    assign n217 = n191 ? sys_r_line[6] : 1'b0;   // memory_op.v(58)
    assign n218 = n191 ? sys_r_line[5] : 1'b1;   // memory_op.v(58)
    assign n219 = n191 ? sys_r_line[4] : 1'b0;   // memory_op.v(58)
    assign n220 = n191 ? sys_r_line[3] : 1'b1;   // memory_op.v(58)
    assign n221 = n191 ? sys_r_line[2] : 1'b0;   // memory_op.v(58)
    assign n222 = n191 ? sys_r_line[1] : 1'b1;   // memory_op.v(58)
    assign n223 = n191 ? sys_r_line[0] : 1'b0;   // memory_op.v(58)
    assign n224 = n189 ? ram_r_line[31] : n192;   // memory_op.v(58)
    assign n225 = n189 ? ram_r_line[30] : n193;   // memory_op.v(58)
    assign n226 = n189 ? ram_r_line[29] : n194;   // memory_op.v(58)
    assign n227 = n189 ? ram_r_line[28] : n195;   // memory_op.v(58)
    assign n228 = n189 ? ram_r_line[27] : n196;   // memory_op.v(58)
    assign n229 = n189 ? ram_r_line[26] : n197;   // memory_op.v(58)
    assign n230 = n189 ? ram_r_line[25] : n198;   // memory_op.v(58)
    assign n231 = n189 ? ram_r_line[24] : n199;   // memory_op.v(58)
    assign n232 = n189 ? ram_r_line[23] : n200;   // memory_op.v(58)
    assign n233 = n189 ? ram_r_line[22] : n201;   // memory_op.v(58)
    assign n234 = n189 ? ram_r_line[21] : n202;   // memory_op.v(58)
    assign n235 = n189 ? ram_r_line[20] : n203;   // memory_op.v(58)
    assign n236 = n189 ? ram_r_line[19] : n204;   // memory_op.v(58)
    assign n237 = n189 ? ram_r_line[18] : n205;   // memory_op.v(58)
    assign n238 = n189 ? ram_r_line[17] : n206;   // memory_op.v(58)
    assign n239 = n189 ? ram_r_line[16] : n207;   // memory_op.v(58)
    assign n240 = n189 ? ram_r_line[15] : n208;   // memory_op.v(58)
    assign n241 = n189 ? ram_r_line[14] : n209;   // memory_op.v(58)
    assign n242 = n189 ? ram_r_line[13] : n210;   // memory_op.v(58)
    assign n243 = n189 ? ram_r_line[12] : n211;   // memory_op.v(58)
    assign n244 = n189 ? ram_r_line[11] : n212;   // memory_op.v(58)
    assign n245 = n189 ? ram_r_line[10] : n213;   // memory_op.v(58)
    assign n246 = n189 ? ram_r_line[9] : n214;   // memory_op.v(58)
    assign n247 = n189 ? ram_r_line[8] : n215;   // memory_op.v(58)
    assign n248 = n189 ? ram_r_line[7] : n216;   // memory_op.v(58)
    assign n249 = n189 ? ram_r_line[6] : n217;   // memory_op.v(58)
    assign n250 = n189 ? ram_r_line[5] : n218;   // memory_op.v(58)
    assign n251 = n189 ? ram_r_line[4] : n219;   // memory_op.v(58)
    assign n252 = n189 ? ram_r_line[3] : n220;   // memory_op.v(58)
    assign n253 = n189 ? ram_r_line[2] : n221;   // memory_op.v(58)
    assign n254 = n189 ? ram_r_line[1] : n222;   // memory_op.v(58)
    assign n255 = n189 ? ram_r_line[0] : n223;   // memory_op.v(58)
    assign n256 = n186 ? r2_inner[31] : n224;   // memory_op.v(58)
    assign n257 = n186 ? r2_inner[30] : n225;   // memory_op.v(58)
    assign n258 = n186 ? r2_inner[29] : n226;   // memory_op.v(58)
    assign n259 = n186 ? r2_inner[28] : n227;   // memory_op.v(58)
    assign n260 = n186 ? r2_inner[27] : n228;   // memory_op.v(58)
    assign n261 = n186 ? r2_inner[26] : n229;   // memory_op.v(58)
    assign n262 = n186 ? r2_inner[25] : n230;   // memory_op.v(58)
    assign n263 = n186 ? r2_inner[24] : n231;   // memory_op.v(58)
    assign n264 = n186 ? r2_inner[23] : n232;   // memory_op.v(58)
    assign n265 = n186 ? r2_inner[22] : n233;   // memory_op.v(58)
    assign n266 = n186 ? r2_inner[21] : n234;   // memory_op.v(58)
    assign n267 = n186 ? r2_inner[20] : n235;   // memory_op.v(58)
    assign n268 = n186 ? r2_inner[19] : n236;   // memory_op.v(58)
    assign n269 = n186 ? r2_inner[18] : n237;   // memory_op.v(58)
    assign n270 = n186 ? r2_inner[17] : n238;   // memory_op.v(58)
    assign n271 = n186 ? r2_inner[16] : n239;   // memory_op.v(58)
    assign n272 = n186 ? r2_inner[15] : n240;   // memory_op.v(58)
    assign n273 = n186 ? r2_inner[14] : n241;   // memory_op.v(58)
    assign n274 = n186 ? r2_inner[13] : n242;   // memory_op.v(58)
    assign n275 = n186 ? r2_inner[12] : n243;   // memory_op.v(58)
    assign n276 = n186 ? r2_inner[11] : n244;   // memory_op.v(58)
    assign n277 = n186 ? r2_inner[10] : n245;   // memory_op.v(58)
    assign n278 = n186 ? r2_inner[9] : n246;   // memory_op.v(58)
    assign n279 = n186 ? r2_inner[8] : n247;   // memory_op.v(58)
    assign n280 = n186 ? r2_inner[7] : n248;   // memory_op.v(58)
    assign n281 = n186 ? r2_inner[6] : n249;   // memory_op.v(58)
    assign n282 = n186 ? r2_inner[5] : n250;   // memory_op.v(58)
    assign n283 = n186 ? r2_inner[4] : n251;   // memory_op.v(58)
    assign n284 = n186 ? r2_inner[3] : n252;   // memory_op.v(58)
    assign n285 = n186 ? r2_inner[2] : n253;   // memory_op.v(58)
    assign n286 = n186 ? r2_inner[1] : n254;   // memory_op.v(58)
    assign n287 = n186 ? r2_inner[0] : n255;   // memory_op.v(58)
    assign n288 = n184 ? r1_inner[31] : n256;   // memory_op.v(58)
    assign n289 = n184 ? r1_inner[30] : n257;   // memory_op.v(58)
    assign n290 = n184 ? r1_inner[29] : n258;   // memory_op.v(58)
    assign n291 = n184 ? r1_inner[28] : n259;   // memory_op.v(58)
    assign n292 = n184 ? r1_inner[27] : n260;   // memory_op.v(58)
    assign n293 = n184 ? r1_inner[26] : n261;   // memory_op.v(58)
    assign n294 = n184 ? r1_inner[25] : n262;   // memory_op.v(58)
    assign n295 = n184 ? r1_inner[24] : n263;   // memory_op.v(58)
    assign n296 = n184 ? r1_inner[23] : n264;   // memory_op.v(58)
    assign n297 = n184 ? r1_inner[22] : n265;   // memory_op.v(58)
    assign n298 = n184 ? r1_inner[21] : n266;   // memory_op.v(58)
    assign n299 = n184 ? r1_inner[20] : n267;   // memory_op.v(58)
    assign n300 = n184 ? r1_inner[19] : n268;   // memory_op.v(58)
    assign n301 = n184 ? r1_inner[18] : n269;   // memory_op.v(58)
    assign n302 = n184 ? r1_inner[17] : n270;   // memory_op.v(58)
    assign n303 = n184 ? r1_inner[16] : n271;   // memory_op.v(58)
    assign n304 = n184 ? r1_inner[15] : n272;   // memory_op.v(58)
    assign n305 = n184 ? r1_inner[14] : n273;   // memory_op.v(58)
    assign n306 = n184 ? r1_inner[13] : n274;   // memory_op.v(58)
    assign n307 = n184 ? r1_inner[12] : n275;   // memory_op.v(58)
    assign n308 = n184 ? r1_inner[11] : n276;   // memory_op.v(58)
    assign n309 = n184 ? r1_inner[10] : n277;   // memory_op.v(58)
    assign n310 = n184 ? r1_inner[9] : n278;   // memory_op.v(58)
    assign n311 = n184 ? r1_inner[8] : n279;   // memory_op.v(58)
    assign n312 = n184 ? r1_inner[7] : n280;   // memory_op.v(58)
    assign n313 = n184 ? r1_inner[6] : n281;   // memory_op.v(58)
    assign n314 = n184 ? r1_inner[5] : n282;   // memory_op.v(58)
    assign n315 = n184 ? r1_inner[4] : n283;   // memory_op.v(58)
    assign n316 = n184 ? r1_inner[3] : n284;   // memory_op.v(58)
    assign n317 = n184 ? r1_inner[2] : n285;   // memory_op.v(58)
    assign n318 = n184 ? r1_inner[1] : n286;   // memory_op.v(58)
    assign n319 = n184 ? r1_inner[0] : n287;   // memory_op.v(58)
    assign m2[31] = n182 ? 1'b0 : n288;   // memory_op.v(58)
    assign m2[30] = n182 ? 1'b0 : n289;   // memory_op.v(58)
    assign m2[29] = n182 ? 1'b0 : n290;   // memory_op.v(58)
    assign m2[28] = n182 ? 1'b0 : n291;   // memory_op.v(58)
    assign m2[27] = n182 ? 1'b0 : n292;   // memory_op.v(58)
    assign m2[26] = n182 ? 1'b0 : n293;   // memory_op.v(58)
    assign m2[25] = n182 ? 1'b0 : n294;   // memory_op.v(58)
    assign m2[24] = n182 ? 1'b0 : n295;   // memory_op.v(58)
    assign m2[23] = n182 ? 1'b0 : n296;   // memory_op.v(58)
    assign m2[22] = n182 ? 1'b0 : n297;   // memory_op.v(58)
    assign m2[21] = n182 ? 1'b0 : n298;   // memory_op.v(58)
    assign m2[20] = n182 ? 1'b0 : n299;   // memory_op.v(58)
    assign m2[19] = n182 ? 1'b0 : n300;   // memory_op.v(58)
    assign m2[18] = n182 ? 1'b0 : n301;   // memory_op.v(58)
    assign m2[17] = n182 ? 1'b0 : n302;   // memory_op.v(58)
    assign m2[16] = n182 ? 1'b0 : n303;   // memory_op.v(58)
    assign m2[15] = n182 ? 1'b0 : n304;   // memory_op.v(58)
    assign m2[14] = n182 ? 1'b0 : n305;   // memory_op.v(58)
    assign m2[13] = n182 ? 1'b0 : n306;   // memory_op.v(58)
    assign m2[12] = n182 ? 1'b0 : n307;   // memory_op.v(58)
    assign m2[11] = n182 ? 1'b0 : n308;   // memory_op.v(58)
    assign m2[10] = n182 ? 1'b0 : n309;   // memory_op.v(58)
    assign m2[9] = n182 ? 1'b0 : n310;   // memory_op.v(58)
    assign m2[8] = n182 ? 1'b0 : n311;   // memory_op.v(58)
    assign m2[7] = n182 ? 1'b0 : n312;   // memory_op.v(58)
    assign m2[6] = n182 ? 1'b0 : n313;   // memory_op.v(58)
    assign m2[5] = n182 ? 1'b0 : n314;   // memory_op.v(58)
    assign m2[4] = n182 ? 1'b0 : n315;   // memory_op.v(58)
    assign m2[3] = n182 ? 1'b0 : n316;   // memory_op.v(58)
    assign m2[2] = n182 ? 1'b0 : n317;   // memory_op.v(58)
    assign m2[1] = n182 ? 1'b0 : n318;   // memory_op.v(58)
    assign m2[0] = n182 ? 1'b0 : n319;   // memory_op.v(58)
    Mux_4u_16u Mux_352 (.sel({r1_op_inner}), .data({m1_select[2], 15'b000011100000000}), 
            .o(n353));   // memory_op.v(73)
    Mux_4u_16u Mux_353 (.sel({r1_op_inner}), .data({m1_select[1], 15'b100000000011100}), 
            .o(n354));   // memory_op.v(73)
    Mux_4u_16u Mux_354 (.sel({r1_op_inner}), .data({m1_select[0], 15'b011100011111110}), 
            .o(n355));   // memory_op.v(73)
    Mux_4u_16u Mux_355 (.sel({r1_op_inner}), .data({sys_w_line[31], sys_w_line[31], 
            r1[31], r1[31], r1[31], sys_w_line[31], sys_w_line[31], 
            sys_w_line[31], sys_w_line[31], sys_w_line[31], sys_w_line[31], 
            sys_w_line[31], sys_w_line[31], sys_w_line[31], sys_w_line[31], 
            sys_w_line[31]}), .o(n356));   // memory_op.v(73)
    Mux_4u_16u Mux_356 (.sel({r1_op_inner}), .data({sys_w_line[30], sys_w_line[30], 
            r1[30], r1[30], r1[30], sys_w_line[30], sys_w_line[30], 
            sys_w_line[30], sys_w_line[30], sys_w_line[30], sys_w_line[30], 
            sys_w_line[30], sys_w_line[30], sys_w_line[30], sys_w_line[30], 
            sys_w_line[30]}), .o(n357));   // memory_op.v(73)
    Mux_4u_16u Mux_357 (.sel({r1_op_inner}), .data({sys_w_line[29], sys_w_line[29], 
            r1[29], r1[29], r1[29], sys_w_line[29], sys_w_line[29], 
            sys_w_line[29], sys_w_line[29], sys_w_line[29], sys_w_line[29], 
            sys_w_line[29], sys_w_line[29], sys_w_line[29], sys_w_line[29], 
            sys_w_line[29]}), .o(n358));   // memory_op.v(73)
    Mux_4u_16u Mux_358 (.sel({r1_op_inner}), .data({sys_w_line[28], sys_w_line[28], 
            r1[28], r1[28], r1[28], sys_w_line[28], sys_w_line[28], 
            sys_w_line[28], sys_w_line[28], sys_w_line[28], sys_w_line[28], 
            sys_w_line[28], sys_w_line[28], sys_w_line[28], sys_w_line[28], 
            sys_w_line[28]}), .o(n359));   // memory_op.v(73)
    Mux_4u_16u Mux_359 (.sel({r1_op_inner}), .data({sys_w_line[27], sys_w_line[27], 
            r1[27], r1[27], r1[27], sys_w_line[27], sys_w_line[27], 
            sys_w_line[27], sys_w_line[27], sys_w_line[27], sys_w_line[27], 
            sys_w_line[27], sys_w_line[27], sys_w_line[27], sys_w_line[27], 
            sys_w_line[27]}), .o(n360));   // memory_op.v(73)
    Mux_4u_16u Mux_360 (.sel({r1_op_inner}), .data({sys_w_line[26], sys_w_line[26], 
            r1[26], r1[26], r1[26], sys_w_line[26], sys_w_line[26], 
            sys_w_line[26], sys_w_line[26], sys_w_line[26], sys_w_line[26], 
            sys_w_line[26], sys_w_line[26], sys_w_line[26], sys_w_line[26], 
            sys_w_line[26]}), .o(n361));   // memory_op.v(73)
    Mux_4u_16u Mux_361 (.sel({r1_op_inner}), .data({sys_w_line[25], sys_w_line[25], 
            r1[25], r1[25], r1[25], sys_w_line[25], sys_w_line[25], 
            sys_w_line[25], sys_w_line[25], sys_w_line[25], sys_w_line[25], 
            sys_w_line[25], sys_w_line[25], sys_w_line[25], sys_w_line[25], 
            sys_w_line[25]}), .o(n362));   // memory_op.v(73)
    Mux_4u_16u Mux_362 (.sel({r1_op_inner}), .data({sys_w_line[24], sys_w_line[24], 
            r1[24], r1[24], r1[24], sys_w_line[24], sys_w_line[24], 
            sys_w_line[24], sys_w_line[24], sys_w_line[24], sys_w_line[24], 
            sys_w_line[24], sys_w_line[24], sys_w_line[24], sys_w_line[24], 
            sys_w_line[24]}), .o(n363));   // memory_op.v(73)
    Mux_4u_16u Mux_363 (.sel({r1_op_inner}), .data({sys_w_line[23], sys_w_line[23], 
            r1[23], r1[23], r1[23], sys_w_line[23], sys_w_line[23], 
            sys_w_line[23], sys_w_line[23], sys_w_line[23], sys_w_line[23], 
            sys_w_line[23], sys_w_line[23], sys_w_line[23], sys_w_line[23], 
            sys_w_line[23]}), .o(n364));   // memory_op.v(73)
    Mux_4u_16u Mux_364 (.sel({r1_op_inner}), .data({sys_w_line[22], sys_w_line[22], 
            r1[22], r1[22], r1[22], sys_w_line[22], sys_w_line[22], 
            sys_w_line[22], sys_w_line[22], sys_w_line[22], sys_w_line[22], 
            sys_w_line[22], sys_w_line[22], sys_w_line[22], sys_w_line[22], 
            sys_w_line[22]}), .o(n365));   // memory_op.v(73)
    Mux_4u_16u Mux_365 (.sel({r1_op_inner}), .data({sys_w_line[21], sys_w_line[21], 
            r1[21], r1[21], r1[21], sys_w_line[21], sys_w_line[21], 
            sys_w_line[21], sys_w_line[21], sys_w_line[21], sys_w_line[21], 
            sys_w_line[21], sys_w_line[21], sys_w_line[21], sys_w_line[21], 
            sys_w_line[21]}), .o(n366));   // memory_op.v(73)
    Mux_4u_16u Mux_366 (.sel({r1_op_inner}), .data({sys_w_line[20], sys_w_line[20], 
            r1[20], r1[20], r1[20], sys_w_line[20], sys_w_line[20], 
            sys_w_line[20], sys_w_line[20], sys_w_line[20], sys_w_line[20], 
            sys_w_line[20], sys_w_line[20], sys_w_line[20], sys_w_line[20], 
            sys_w_line[20]}), .o(n367));   // memory_op.v(73)
    Mux_4u_16u Mux_367 (.sel({r1_op_inner}), .data({sys_w_line[19], sys_w_line[19], 
            r1[19], r1[19], r1[19], sys_w_line[19], sys_w_line[19], 
            sys_w_line[19], sys_w_line[19], sys_w_line[19], sys_w_line[19], 
            sys_w_line[19], sys_w_line[19], sys_w_line[19], sys_w_line[19], 
            sys_w_line[19]}), .o(n368));   // memory_op.v(73)
    Mux_4u_16u Mux_368 (.sel({r1_op_inner}), .data({sys_w_line[18], sys_w_line[18], 
            r1[18], r1[18], r1[18], sys_w_line[18], sys_w_line[18], 
            sys_w_line[18], sys_w_line[18], sys_w_line[18], sys_w_line[18], 
            sys_w_line[18], sys_w_line[18], sys_w_line[18], sys_w_line[18], 
            sys_w_line[18]}), .o(n369));   // memory_op.v(73)
    Mux_4u_16u Mux_369 (.sel({r1_op_inner}), .data({sys_w_line[17], sys_w_line[17], 
            r1[17], r1[17], r1[17], sys_w_line[17], sys_w_line[17], 
            sys_w_line[17], sys_w_line[17], sys_w_line[17], sys_w_line[17], 
            sys_w_line[17], sys_w_line[17], sys_w_line[17], sys_w_line[17], 
            sys_w_line[17]}), .o(n370));   // memory_op.v(73)
    Mux_4u_16u Mux_370 (.sel({r1_op_inner}), .data({sys_w_line[16], sys_w_line[16], 
            r1[16], r1[16], r1[16], sys_w_line[16], sys_w_line[16], 
            sys_w_line[16], sys_w_line[16], sys_w_line[16], sys_w_line[16], 
            sys_w_line[16], sys_w_line[16], sys_w_line[16], sys_w_line[16], 
            sys_w_line[16]}), .o(n371));   // memory_op.v(73)
    Mux_4u_16u Mux_371 (.sel({r1_op_inner}), .data({sys_w_line[15], sys_w_line[15], 
            r1[15], r1[15], r1[15], sys_w_line[15], sys_w_line[15], 
            sys_w_line[15], sys_w_line[15], sys_w_line[15], sys_w_line[15], 
            sys_w_line[15], sys_w_line[15], sys_w_line[15], sys_w_line[15], 
            sys_w_line[15]}), .o(n372));   // memory_op.v(73)
    Mux_4u_16u Mux_372 (.sel({r1_op_inner}), .data({sys_w_line[14], sys_w_line[14], 
            r1[14], r1[14], r1[14], sys_w_line[14], sys_w_line[14], 
            sys_w_line[14], sys_w_line[14], sys_w_line[14], sys_w_line[14], 
            sys_w_line[14], sys_w_line[14], sys_w_line[14], sys_w_line[14], 
            sys_w_line[14]}), .o(n373));   // memory_op.v(73)
    Mux_4u_16u Mux_373 (.sel({r1_op_inner}), .data({sys_w_line[13], sys_w_line[13], 
            r1[13], r1[13], r1[13], sys_w_line[13], sys_w_line[13], 
            sys_w_line[13], sys_w_line[13], sys_w_line[13], sys_w_line[13], 
            sys_w_line[13], sys_w_line[13], sys_w_line[13], sys_w_line[13], 
            sys_w_line[13]}), .o(n374));   // memory_op.v(73)
    Mux_4u_16u Mux_374 (.sel({r1_op_inner}), .data({sys_w_line[12], sys_w_line[12], 
            r1[12], r1[12], r1[12], sys_w_line[12], sys_w_line[12], 
            sys_w_line[12], sys_w_line[12], sys_w_line[12], sys_w_line[12], 
            sys_w_line[12], sys_w_line[12], sys_w_line[12], sys_w_line[12], 
            sys_w_line[12]}), .o(n375));   // memory_op.v(73)
    Mux_4u_16u Mux_375 (.sel({r1_op_inner}), .data({sys_w_line[11], sys_w_line[11], 
            r1[11], r1[11], r1[11], sys_w_line[11], sys_w_line[11], 
            sys_w_line[11], sys_w_line[11], sys_w_line[11], sys_w_line[11], 
            sys_w_line[11], sys_w_line[11], sys_w_line[11], sys_w_line[11], 
            sys_w_line[11]}), .o(n376));   // memory_op.v(73)
    Mux_4u_16u Mux_376 (.sel({r1_op_inner}), .data({sys_w_line[10], sys_w_line[10], 
            r1[10], r1[10], r1[10], sys_w_line[10], sys_w_line[10], 
            sys_w_line[10], sys_w_line[10], sys_w_line[10], sys_w_line[10], 
            sys_w_line[10], sys_w_line[10], sys_w_line[10], sys_w_line[10], 
            sys_w_line[10]}), .o(n377));   // memory_op.v(73)
    Mux_4u_16u Mux_377 (.sel({r1_op_inner}), .data({sys_w_line[9], sys_w_line[9], 
            r1[9], r1[9], r1[9], sys_w_line[9], sys_w_line[9], sys_w_line[9], 
            sys_w_line[9], sys_w_line[9], sys_w_line[9], sys_w_line[9], 
            sys_w_line[9], sys_w_line[9], sys_w_line[9], sys_w_line[9]}), 
            .o(n378));   // memory_op.v(73)
    Mux_4u_16u Mux_378 (.sel({r1_op_inner}), .data({sys_w_line[8], sys_w_line[8], 
            r1[8], r1[8], r1[8], sys_w_line[8], sys_w_line[8], sys_w_line[8], 
            sys_w_line[8], sys_w_line[8], sys_w_line[8], sys_w_line[8], 
            sys_w_line[8], sys_w_line[8], sys_w_line[8], sys_w_line[8]}), 
            .o(n379));   // memory_op.v(73)
    Mux_4u_16u Mux_379 (.sel({r1_op_inner}), .data({sys_w_line[7], sys_w_line[7], 
            r1[7], r1[7], r1[7], sys_w_line[7], sys_w_line[7], sys_w_line[7], 
            sys_w_line[7], sys_w_line[7], sys_w_line[7], sys_w_line[7], 
            sys_w_line[7], sys_w_line[7], sys_w_line[7], sys_w_line[7]}), 
            .o(n380));   // memory_op.v(73)
    Mux_4u_16u Mux_380 (.sel({r1_op_inner}), .data({sys_w_line[6], sys_w_line[6], 
            r1[6], r1[6], r1[6], sys_w_line[6], sys_w_line[6], sys_w_line[6], 
            sys_w_line[6], sys_w_line[6], sys_w_line[6], sys_w_line[6], 
            sys_w_line[6], sys_w_line[6], sys_w_line[6], sys_w_line[6]}), 
            .o(n381));   // memory_op.v(73)
    Mux_4u_16u Mux_381 (.sel({r1_op_inner}), .data({sys_w_line[5], sys_w_line[5], 
            r1[5], r1[5], r1[5], sys_w_line[5], sys_w_line[5], sys_w_line[5], 
            sys_w_line[5], sys_w_line[5], sys_w_line[5], sys_w_line[5], 
            sys_w_line[5], sys_w_line[5], sys_w_line[5], sys_w_line[5]}), 
            .o(n382));   // memory_op.v(73)
    Mux_4u_16u Mux_382 (.sel({r1_op_inner}), .data({sys_w_line[4], sys_w_line[4], 
            r1[4], r1[4], r1[4], sys_w_line[4], sys_w_line[4], sys_w_line[4], 
            sys_w_line[4], sys_w_line[4], sys_w_line[4], sys_w_line[4], 
            sys_w_line[4], sys_w_line[4], sys_w_line[4], sys_w_line[4]}), 
            .o(n383));   // memory_op.v(73)
    Mux_4u_16u Mux_383 (.sel({r1_op_inner}), .data({sys_w_line[3], sys_w_line[3], 
            r1[3], r1[3], r1[3], sys_w_line[3], sys_w_line[3], sys_w_line[3], 
            sys_w_line[3], sys_w_line[3], sys_w_line[3], sys_w_line[3], 
            sys_w_line[3], sys_w_line[3], sys_w_line[3], sys_w_line[3]}), 
            .o(n384));   // memory_op.v(73)
    Mux_4u_16u Mux_384 (.sel({r1_op_inner}), .data({sys_w_line[2], sys_w_line[2], 
            r1[2], r1[2], r1[2], sys_w_line[2], sys_w_line[2], sys_w_line[2], 
            sys_w_line[2], sys_w_line[2], sys_w_line[2], sys_w_line[2], 
            sys_w_line[2], sys_w_line[2], sys_w_line[2], sys_w_line[2]}), 
            .o(n385));   // memory_op.v(73)
    Mux_4u_16u Mux_385 (.sel({r1_op_inner}), .data({sys_w_line[1], sys_w_line[1], 
            r1[1], r1[1], r1[1], sys_w_line[1], sys_w_line[1], sys_w_line[1], 
            sys_w_line[1], sys_w_line[1], sys_w_line[1], sys_w_line[1], 
            sys_w_line[1], sys_w_line[1], sys_w_line[1], sys_w_line[1]}), 
            .o(n386));   // memory_op.v(73)
    Mux_4u_16u Mux_386 (.sel({r1_op_inner}), .data({sys_w_line[0], sys_w_line[0], 
            r1[0], r1[0], r1[0], sys_w_line[0], sys_w_line[0], sys_w_line[0], 
            sys_w_line[0], sys_w_line[0], sys_w_line[0], sys_w_line[0], 
            sys_w_line[0], sys_w_line[0], sys_w_line[0], sys_w_line[0]}), 
            .o(n387));   // memory_op.v(73)
    Mux_4u_16u Mux_387 (.sel({r1_op_inner}), .data({sys_w_addr[31], sys_w_addr[31], 
            r2[31], a2[31], a1[31], sys_w_addr[31], sys_w_addr[31], 
            sys_w_addr[31], sys_w_addr[31], sys_w_addr[31], sys_w_addr[31], 
            sys_w_addr[31], sys_w_addr[31], sys_w_addr[31], sys_w_addr[31], 
            sys_w_addr[31]}), .o(n388));   // memory_op.v(73)
    Mux_4u_16u Mux_388 (.sel({r1_op_inner}), .data({sys_w_addr[30], sys_w_addr[30], 
            r2[30], a2[30], a1[30], sys_w_addr[30], sys_w_addr[30], 
            sys_w_addr[30], sys_w_addr[30], sys_w_addr[30], sys_w_addr[30], 
            sys_w_addr[30], sys_w_addr[30], sys_w_addr[30], sys_w_addr[30], 
            sys_w_addr[30]}), .o(n389));   // memory_op.v(73)
    Mux_4u_16u Mux_389 (.sel({r1_op_inner}), .data({sys_w_addr[29], sys_w_addr[29], 
            r2[29], a2[29], a1[29], sys_w_addr[29], sys_w_addr[29], 
            sys_w_addr[29], sys_w_addr[29], sys_w_addr[29], sys_w_addr[29], 
            sys_w_addr[29], sys_w_addr[29], sys_w_addr[29], sys_w_addr[29], 
            sys_w_addr[29]}), .o(n390));   // memory_op.v(73)
    Mux_4u_16u Mux_390 (.sel({r1_op_inner}), .data({sys_w_addr[28], sys_w_addr[28], 
            r2[28], a2[28], a1[28], sys_w_addr[28], sys_w_addr[28], 
            sys_w_addr[28], sys_w_addr[28], sys_w_addr[28], sys_w_addr[28], 
            sys_w_addr[28], sys_w_addr[28], sys_w_addr[28], sys_w_addr[28], 
            sys_w_addr[28]}), .o(n391));   // memory_op.v(73)
    Mux_4u_16u Mux_391 (.sel({r1_op_inner}), .data({sys_w_addr[27], sys_w_addr[27], 
            r2[27], a2[27], a1[27], sys_w_addr[27], sys_w_addr[27], 
            sys_w_addr[27], sys_w_addr[27], sys_w_addr[27], sys_w_addr[27], 
            sys_w_addr[27], sys_w_addr[27], sys_w_addr[27], sys_w_addr[27], 
            sys_w_addr[27]}), .o(n392));   // memory_op.v(73)
    Mux_4u_16u Mux_392 (.sel({r1_op_inner}), .data({sys_w_addr[26], sys_w_addr[26], 
            r2[26], a2[26], a1[26], sys_w_addr[26], sys_w_addr[26], 
            sys_w_addr[26], sys_w_addr[26], sys_w_addr[26], sys_w_addr[26], 
            sys_w_addr[26], sys_w_addr[26], sys_w_addr[26], sys_w_addr[26], 
            sys_w_addr[26]}), .o(n393));   // memory_op.v(73)
    Mux_4u_16u Mux_393 (.sel({r1_op_inner}), .data({sys_w_addr[25], sys_w_addr[25], 
            r2[25], a2[25], a1[25], sys_w_addr[25], sys_w_addr[25], 
            sys_w_addr[25], sys_w_addr[25], sys_w_addr[25], sys_w_addr[25], 
            sys_w_addr[25], sys_w_addr[25], sys_w_addr[25], sys_w_addr[25], 
            sys_w_addr[25]}), .o(n394));   // memory_op.v(73)
    Mux_4u_16u Mux_394 (.sel({r1_op_inner}), .data({sys_w_addr[24], sys_w_addr[24], 
            r2[24], a2[24], a1[24], sys_w_addr[24], sys_w_addr[24], 
            sys_w_addr[24], sys_w_addr[24], sys_w_addr[24], sys_w_addr[24], 
            sys_w_addr[24], sys_w_addr[24], sys_w_addr[24], sys_w_addr[24], 
            sys_w_addr[24]}), .o(n395));   // memory_op.v(73)
    Mux_4u_16u Mux_395 (.sel({r1_op_inner}), .data({sys_w_addr[23], sys_w_addr[23], 
            r2[23], a2[23], a1[23], sys_w_addr[23], sys_w_addr[23], 
            sys_w_addr[23], sys_w_addr[23], sys_w_addr[23], sys_w_addr[23], 
            sys_w_addr[23], sys_w_addr[23], sys_w_addr[23], sys_w_addr[23], 
            sys_w_addr[23]}), .o(n396));   // memory_op.v(73)
    Mux_4u_16u Mux_396 (.sel({r1_op_inner}), .data({sys_w_addr[22], sys_w_addr[22], 
            r2[22], a2[22], a1[22], sys_w_addr[22], sys_w_addr[22], 
            sys_w_addr[22], sys_w_addr[22], sys_w_addr[22], sys_w_addr[22], 
            sys_w_addr[22], sys_w_addr[22], sys_w_addr[22], sys_w_addr[22], 
            sys_w_addr[22]}), .o(n397));   // memory_op.v(73)
    Mux_4u_16u Mux_397 (.sel({r1_op_inner}), .data({sys_w_addr[21], sys_w_addr[21], 
            r2[21], a2[21], a1[21], sys_w_addr[21], sys_w_addr[21], 
            sys_w_addr[21], sys_w_addr[21], sys_w_addr[21], sys_w_addr[21], 
            sys_w_addr[21], sys_w_addr[21], sys_w_addr[21], sys_w_addr[21], 
            sys_w_addr[21]}), .o(n398));   // memory_op.v(73)
    Mux_4u_16u Mux_398 (.sel({r1_op_inner}), .data({sys_w_addr[20], sys_w_addr[20], 
            r2[20], a2[20], a1[20], sys_w_addr[20], sys_w_addr[20], 
            sys_w_addr[20], sys_w_addr[20], sys_w_addr[20], sys_w_addr[20], 
            sys_w_addr[20], sys_w_addr[20], sys_w_addr[20], sys_w_addr[20], 
            sys_w_addr[20]}), .o(n399));   // memory_op.v(73)
    Mux_4u_16u Mux_399 (.sel({r1_op_inner}), .data({sys_w_addr[19], sys_w_addr[19], 
            r2[19], a2[19], a1[19], sys_w_addr[19], sys_w_addr[19], 
            sys_w_addr[19], sys_w_addr[19], sys_w_addr[19], sys_w_addr[19], 
            sys_w_addr[19], sys_w_addr[19], sys_w_addr[19], sys_w_addr[19], 
            sys_w_addr[19]}), .o(n400));   // memory_op.v(73)
    Mux_4u_16u Mux_400 (.sel({r1_op_inner}), .data({sys_w_addr[18], sys_w_addr[18], 
            r2[18], a2[18], a1[18], sys_w_addr[18], sys_w_addr[18], 
            sys_w_addr[18], sys_w_addr[18], sys_w_addr[18], sys_w_addr[18], 
            sys_w_addr[18], sys_w_addr[18], sys_w_addr[18], sys_w_addr[18], 
            sys_w_addr[18]}), .o(n401));   // memory_op.v(73)
    Mux_4u_16u Mux_401 (.sel({r1_op_inner}), .data({sys_w_addr[17], sys_w_addr[17], 
            r2[17], a2[17], a1[17], sys_w_addr[17], sys_w_addr[17], 
            sys_w_addr[17], sys_w_addr[17], sys_w_addr[17], sys_w_addr[17], 
            sys_w_addr[17], sys_w_addr[17], sys_w_addr[17], sys_w_addr[17], 
            sys_w_addr[17]}), .o(n402));   // memory_op.v(73)
    Mux_4u_16u Mux_402 (.sel({r1_op_inner}), .data({sys_w_addr[16], sys_w_addr[16], 
            r2[16], a2[16], a1[16], sys_w_addr[16], sys_w_addr[16], 
            sys_w_addr[16], sys_w_addr[16], sys_w_addr[16], sys_w_addr[16], 
            sys_w_addr[16], sys_w_addr[16], sys_w_addr[16], sys_w_addr[16], 
            sys_w_addr[16]}), .o(n403));   // memory_op.v(73)
    Mux_4u_16u Mux_403 (.sel({r1_op_inner}), .data({sys_w_addr[15], sys_w_addr[15], 
            r2[15], a2[15], a1[15], sys_w_addr[15], sys_w_addr[15], 
            sys_w_addr[15], sys_w_addr[15], sys_w_addr[15], sys_w_addr[15], 
            sys_w_addr[15], sys_w_addr[15], sys_w_addr[15], sys_w_addr[15], 
            sys_w_addr[15]}), .o(n404));   // memory_op.v(73)
    Mux_4u_16u Mux_404 (.sel({r1_op_inner}), .data({sys_w_addr[14], sys_w_addr[14], 
            r2[14], a2[14], a1[14], sys_w_addr[14], sys_w_addr[14], 
            sys_w_addr[14], sys_w_addr[14], sys_w_addr[14], sys_w_addr[14], 
            sys_w_addr[14], sys_w_addr[14], sys_w_addr[14], sys_w_addr[14], 
            sys_w_addr[14]}), .o(n405));   // memory_op.v(73)
    Mux_4u_16u Mux_405 (.sel({r1_op_inner}), .data({sys_w_addr[13], sys_w_addr[13], 
            r2[13], a2[13], a1[13], sys_w_addr[13], sys_w_addr[13], 
            sys_w_addr[13], sys_w_addr[13], sys_w_addr[13], sys_w_addr[13], 
            sys_w_addr[13], sys_w_addr[13], sys_w_addr[13], sys_w_addr[13], 
            sys_w_addr[13]}), .o(n406));   // memory_op.v(73)
    Mux_4u_16u Mux_406 (.sel({r1_op_inner}), .data({sys_w_addr[12], sys_w_addr[12], 
            r2[12], a2[12], a1[12], sys_w_addr[12], sys_w_addr[12], 
            sys_w_addr[12], sys_w_addr[12], sys_w_addr[12], sys_w_addr[12], 
            sys_w_addr[12], sys_w_addr[12], sys_w_addr[12], sys_w_addr[12], 
            sys_w_addr[12]}), .o(n407));   // memory_op.v(73)
    Mux_4u_16u Mux_407 (.sel({r1_op_inner}), .data({sys_w_addr[11], sys_w_addr[11], 
            r2[11], a2[11], a1[11], sys_w_addr[11], sys_w_addr[11], 
            sys_w_addr[11], sys_w_addr[11], sys_w_addr[11], sys_w_addr[11], 
            sys_w_addr[11], sys_w_addr[11], sys_w_addr[11], sys_w_addr[11], 
            sys_w_addr[11]}), .o(n408));   // memory_op.v(73)
    Mux_4u_16u Mux_408 (.sel({r1_op_inner}), .data({sys_w_addr[10], sys_w_addr[10], 
            r2[10], a2[10], a1[10], sys_w_addr[10], sys_w_addr[10], 
            sys_w_addr[10], sys_w_addr[10], sys_w_addr[10], sys_w_addr[10], 
            sys_w_addr[10], sys_w_addr[10], sys_w_addr[10], sys_w_addr[10], 
            sys_w_addr[10]}), .o(n409));   // memory_op.v(73)
    Mux_4u_16u Mux_409 (.sel({r1_op_inner}), .data({sys_w_addr[9], sys_w_addr[9], 
            r2[9], a2[9], a1[9], sys_w_addr[9], sys_w_addr[9], sys_w_addr[9], 
            sys_w_addr[9], sys_w_addr[9], sys_w_addr[9], sys_w_addr[9], 
            sys_w_addr[9], sys_w_addr[9], sys_w_addr[9], sys_w_addr[9]}), 
            .o(n410));   // memory_op.v(73)
    Mux_4u_16u Mux_410 (.sel({r1_op_inner}), .data({sys_w_addr[8], sys_w_addr[8], 
            r2[8], a2[8], a1[8], sys_w_addr[8], sys_w_addr[8], sys_w_addr[8], 
            sys_w_addr[8], sys_w_addr[8], sys_w_addr[8], sys_w_addr[8], 
            sys_w_addr[8], sys_w_addr[8], sys_w_addr[8], sys_w_addr[8]}), 
            .o(n411));   // memory_op.v(73)
    Mux_4u_16u Mux_411 (.sel({r1_op_inner}), .data({sys_w_addr[7], sys_w_addr[7], 
            r2[7], a2[7], a1[7], sys_w_addr[7], sys_w_addr[7], sys_w_addr[7], 
            sys_w_addr[7], sys_w_addr[7], sys_w_addr[7], sys_w_addr[7], 
            sys_w_addr[7], sys_w_addr[7], sys_w_addr[7], sys_w_addr[7]}), 
            .o(n412));   // memory_op.v(73)
    Mux_4u_16u Mux_412 (.sel({r1_op_inner}), .data({sys_w_addr[6], sys_w_addr[6], 
            r2[6], a2[6], a1[6], sys_w_addr[6], sys_w_addr[6], sys_w_addr[6], 
            sys_w_addr[6], sys_w_addr[6], sys_w_addr[6], sys_w_addr[6], 
            sys_w_addr[6], sys_w_addr[6], sys_w_addr[6], sys_w_addr[6]}), 
            .o(n413));   // memory_op.v(73)
    Mux_4u_16u Mux_413 (.sel({r1_op_inner}), .data({sys_w_addr[5], sys_w_addr[5], 
            r2[5], a2[5], a1[5], sys_w_addr[5], sys_w_addr[5], sys_w_addr[5], 
            sys_w_addr[5], sys_w_addr[5], sys_w_addr[5], sys_w_addr[5], 
            sys_w_addr[5], sys_w_addr[5], sys_w_addr[5], sys_w_addr[5]}), 
            .o(n414));   // memory_op.v(73)
    Mux_4u_16u Mux_414 (.sel({r1_op_inner}), .data({sys_w_addr[4], sys_w_addr[4], 
            r2[4], a2[4], a1[4], sys_w_addr[4], sys_w_addr[4], sys_w_addr[4], 
            sys_w_addr[4], sys_w_addr[4], sys_w_addr[4], sys_w_addr[4], 
            sys_w_addr[4], sys_w_addr[4], sys_w_addr[4], sys_w_addr[4]}), 
            .o(n415));   // memory_op.v(73)
    Mux_4u_16u Mux_415 (.sel({r1_op_inner}), .data({sys_w_addr[3], sys_w_addr[3], 
            r2[3], a2[3], a1[3], sys_w_addr[3], sys_w_addr[3], sys_w_addr[3], 
            sys_w_addr[3], sys_w_addr[3], sys_w_addr[3], sys_w_addr[3], 
            sys_w_addr[3], sys_w_addr[3], sys_w_addr[3], sys_w_addr[3]}), 
            .o(n416));   // memory_op.v(73)
    Mux_4u_16u Mux_416 (.sel({r1_op_inner}), .data({sys_w_addr[2], sys_w_addr[2], 
            r2[2], a2[2], a1[2], sys_w_addr[2], sys_w_addr[2], sys_w_addr[2], 
            sys_w_addr[2], sys_w_addr[2], sys_w_addr[2], sys_w_addr[2], 
            sys_w_addr[2], sys_w_addr[2], sys_w_addr[2], sys_w_addr[2]}), 
            .o(n417));   // memory_op.v(73)
    Mux_4u_16u Mux_417 (.sel({r1_op_inner}), .data({sys_w_addr[1], sys_w_addr[1], 
            r2[1], a2[1], a1[1], sys_w_addr[1], sys_w_addr[1], sys_w_addr[1], 
            sys_w_addr[1], sys_w_addr[1], sys_w_addr[1], sys_w_addr[1], 
            sys_w_addr[1], sys_w_addr[1], sys_w_addr[1], sys_w_addr[1]}), 
            .o(n418));   // memory_op.v(73)
    Mux_4u_16u Mux_418 (.sel({r1_op_inner}), .data({sys_w_addr[0], sys_w_addr[0], 
            r2[0], a2[0], a1[0], sys_w_addr[0], sys_w_addr[0], sys_w_addr[0], 
            sys_w_addr[0], sys_w_addr[0], sys_w_addr[0], sys_w_addr[0], 
            sys_w_addr[0], sys_w_addr[0], sys_w_addr[0], sys_w_addr[0]}), 
            .o(n419));   // memory_op.v(73)
    Mux_4u_16u Mux_419 (.sel({r1_op_inner}), .data({16'b0011100000000000}), 
            .o(n420));   // memory_op.v(73)
    Mux_4u_16u Mux_420 (.sel({r1_op_inner}), .data({sys_r_addr[31], sys_r_addr[31], 
            sys_r_addr[31], sys_r_addr[31], sys_r_addr[31], r2[31], 
            a2[31], a1[31], sys_r_addr[31], sys_r_addr[31], sys_r_addr[31], 
            sys_r_addr[31], sys_r_addr[31], sys_r_addr[31], sys_r_addr[31], 
            sys_r_addr[31]}), .o(n421));   // memory_op.v(73)
    Mux_4u_16u Mux_421 (.sel({r1_op_inner}), .data({sys_r_addr[30], sys_r_addr[30], 
            sys_r_addr[30], sys_r_addr[30], sys_r_addr[30], r2[30], 
            a2[30], a1[30], sys_r_addr[30], sys_r_addr[30], sys_r_addr[30], 
            sys_r_addr[30], sys_r_addr[30], sys_r_addr[30], sys_r_addr[30], 
            sys_r_addr[30]}), .o(n422));   // memory_op.v(73)
    Mux_4u_16u Mux_422 (.sel({r1_op_inner}), .data({sys_r_addr[29], sys_r_addr[29], 
            sys_r_addr[29], sys_r_addr[29], sys_r_addr[29], r2[29], 
            a2[29], a1[29], sys_r_addr[29], sys_r_addr[29], sys_r_addr[29], 
            sys_r_addr[29], sys_r_addr[29], sys_r_addr[29], sys_r_addr[29], 
            sys_r_addr[29]}), .o(n423));   // memory_op.v(73)
    Mux_4u_16u Mux_423 (.sel({r1_op_inner}), .data({sys_r_addr[28], sys_r_addr[28], 
            sys_r_addr[28], sys_r_addr[28], sys_r_addr[28], r2[28], 
            a2[28], a1[28], sys_r_addr[28], sys_r_addr[28], sys_r_addr[28], 
            sys_r_addr[28], sys_r_addr[28], sys_r_addr[28], sys_r_addr[28], 
            sys_r_addr[28]}), .o(n424));   // memory_op.v(73)
    Mux_4u_16u Mux_424 (.sel({r1_op_inner}), .data({sys_r_addr[27], sys_r_addr[27], 
            sys_r_addr[27], sys_r_addr[27], sys_r_addr[27], r2[27], 
            a2[27], a1[27], sys_r_addr[27], sys_r_addr[27], sys_r_addr[27], 
            sys_r_addr[27], sys_r_addr[27], sys_r_addr[27], sys_r_addr[27], 
            sys_r_addr[27]}), .o(n425));   // memory_op.v(73)
    Mux_4u_16u Mux_425 (.sel({r1_op_inner}), .data({sys_r_addr[26], sys_r_addr[26], 
            sys_r_addr[26], sys_r_addr[26], sys_r_addr[26], r2[26], 
            a2[26], a1[26], sys_r_addr[26], sys_r_addr[26], sys_r_addr[26], 
            sys_r_addr[26], sys_r_addr[26], sys_r_addr[26], sys_r_addr[26], 
            sys_r_addr[26]}), .o(n426));   // memory_op.v(73)
    Mux_4u_16u Mux_426 (.sel({r1_op_inner}), .data({sys_r_addr[25], sys_r_addr[25], 
            sys_r_addr[25], sys_r_addr[25], sys_r_addr[25], r2[25], 
            a2[25], a1[25], sys_r_addr[25], sys_r_addr[25], sys_r_addr[25], 
            sys_r_addr[25], sys_r_addr[25], sys_r_addr[25], sys_r_addr[25], 
            sys_r_addr[25]}), .o(n427));   // memory_op.v(73)
    Mux_4u_16u Mux_427 (.sel({r1_op_inner}), .data({sys_r_addr[24], sys_r_addr[24], 
            sys_r_addr[24], sys_r_addr[24], sys_r_addr[24], r2[24], 
            a2[24], a1[24], sys_r_addr[24], sys_r_addr[24], sys_r_addr[24], 
            sys_r_addr[24], sys_r_addr[24], sys_r_addr[24], sys_r_addr[24], 
            sys_r_addr[24]}), .o(n428));   // memory_op.v(73)
    Mux_4u_16u Mux_428 (.sel({r1_op_inner}), .data({sys_r_addr[23], sys_r_addr[23], 
            sys_r_addr[23], sys_r_addr[23], sys_r_addr[23], r2[23], 
            a2[23], a1[23], sys_r_addr[23], sys_r_addr[23], sys_r_addr[23], 
            sys_r_addr[23], sys_r_addr[23], sys_r_addr[23], sys_r_addr[23], 
            sys_r_addr[23]}), .o(n429));   // memory_op.v(73)
    Mux_4u_16u Mux_429 (.sel({r1_op_inner}), .data({sys_r_addr[22], sys_r_addr[22], 
            sys_r_addr[22], sys_r_addr[22], sys_r_addr[22], r2[22], 
            a2[22], a1[22], sys_r_addr[22], sys_r_addr[22], sys_r_addr[22], 
            sys_r_addr[22], sys_r_addr[22], sys_r_addr[22], sys_r_addr[22], 
            sys_r_addr[22]}), .o(n430));   // memory_op.v(73)
    Mux_4u_16u Mux_430 (.sel({r1_op_inner}), .data({sys_r_addr[21], sys_r_addr[21], 
            sys_r_addr[21], sys_r_addr[21], sys_r_addr[21], r2[21], 
            a2[21], a1[21], sys_r_addr[21], sys_r_addr[21], sys_r_addr[21], 
            sys_r_addr[21], sys_r_addr[21], sys_r_addr[21], sys_r_addr[21], 
            sys_r_addr[21]}), .o(n431));   // memory_op.v(73)
    Mux_4u_16u Mux_431 (.sel({r1_op_inner}), .data({sys_r_addr[20], sys_r_addr[20], 
            sys_r_addr[20], sys_r_addr[20], sys_r_addr[20], r2[20], 
            a2[20], a1[20], sys_r_addr[20], sys_r_addr[20], sys_r_addr[20], 
            sys_r_addr[20], sys_r_addr[20], sys_r_addr[20], sys_r_addr[20], 
            sys_r_addr[20]}), .o(n432));   // memory_op.v(73)
    Mux_4u_16u Mux_432 (.sel({r1_op_inner}), .data({sys_r_addr[19], sys_r_addr[19], 
            sys_r_addr[19], sys_r_addr[19], sys_r_addr[19], r2[19], 
            a2[19], a1[19], sys_r_addr[19], sys_r_addr[19], sys_r_addr[19], 
            sys_r_addr[19], sys_r_addr[19], sys_r_addr[19], sys_r_addr[19], 
            sys_r_addr[19]}), .o(n433));   // memory_op.v(73)
    Mux_4u_16u Mux_433 (.sel({r1_op_inner}), .data({sys_r_addr[18], sys_r_addr[18], 
            sys_r_addr[18], sys_r_addr[18], sys_r_addr[18], r2[18], 
            a2[18], a1[18], sys_r_addr[18], sys_r_addr[18], sys_r_addr[18], 
            sys_r_addr[18], sys_r_addr[18], sys_r_addr[18], sys_r_addr[18], 
            sys_r_addr[18]}), .o(n434));   // memory_op.v(73)
    Mux_4u_16u Mux_434 (.sel({r1_op_inner}), .data({sys_r_addr[17], sys_r_addr[17], 
            sys_r_addr[17], sys_r_addr[17], sys_r_addr[17], r2[17], 
            a2[17], a1[17], sys_r_addr[17], sys_r_addr[17], sys_r_addr[17], 
            sys_r_addr[17], sys_r_addr[17], sys_r_addr[17], sys_r_addr[17], 
            sys_r_addr[17]}), .o(n435));   // memory_op.v(73)
    Mux_4u_16u Mux_435 (.sel({r1_op_inner}), .data({sys_r_addr[16], sys_r_addr[16], 
            sys_r_addr[16], sys_r_addr[16], sys_r_addr[16], r2[16], 
            a2[16], a1[16], sys_r_addr[16], sys_r_addr[16], sys_r_addr[16], 
            sys_r_addr[16], sys_r_addr[16], sys_r_addr[16], sys_r_addr[16], 
            sys_r_addr[16]}), .o(n436));   // memory_op.v(73)
    Mux_4u_16u Mux_436 (.sel({r1_op_inner}), .data({sys_r_addr[15], sys_r_addr[15], 
            sys_r_addr[15], sys_r_addr[15], sys_r_addr[15], r2[15], 
            a2[15], a1[15], sys_r_addr[15], sys_r_addr[15], sys_r_addr[15], 
            sys_r_addr[15], sys_r_addr[15], sys_r_addr[15], sys_r_addr[15], 
            sys_r_addr[15]}), .o(n437));   // memory_op.v(73)
    Mux_4u_16u Mux_437 (.sel({r1_op_inner}), .data({sys_r_addr[14], sys_r_addr[14], 
            sys_r_addr[14], sys_r_addr[14], sys_r_addr[14], r2[14], 
            a2[14], a1[14], sys_r_addr[14], sys_r_addr[14], sys_r_addr[14], 
            sys_r_addr[14], sys_r_addr[14], sys_r_addr[14], sys_r_addr[14], 
            sys_r_addr[14]}), .o(n438));   // memory_op.v(73)
    Mux_4u_16u Mux_438 (.sel({r1_op_inner}), .data({sys_r_addr[13], sys_r_addr[13], 
            sys_r_addr[13], sys_r_addr[13], sys_r_addr[13], r2[13], 
            a2[13], a1[13], sys_r_addr[13], sys_r_addr[13], sys_r_addr[13], 
            sys_r_addr[13], sys_r_addr[13], sys_r_addr[13], sys_r_addr[13], 
            sys_r_addr[13]}), .o(n439));   // memory_op.v(73)
    Mux_4u_16u Mux_439 (.sel({r1_op_inner}), .data({sys_r_addr[12], sys_r_addr[12], 
            sys_r_addr[12], sys_r_addr[12], sys_r_addr[12], r2[12], 
            a2[12], a1[12], sys_r_addr[12], sys_r_addr[12], sys_r_addr[12], 
            sys_r_addr[12], sys_r_addr[12], sys_r_addr[12], sys_r_addr[12], 
            sys_r_addr[12]}), .o(n440));   // memory_op.v(73)
    Mux_4u_16u Mux_440 (.sel({r1_op_inner}), .data({sys_r_addr[11], sys_r_addr[11], 
            sys_r_addr[11], sys_r_addr[11], sys_r_addr[11], r2[11], 
            a2[11], a1[11], sys_r_addr[11], sys_r_addr[11], sys_r_addr[11], 
            sys_r_addr[11], sys_r_addr[11], sys_r_addr[11], sys_r_addr[11], 
            sys_r_addr[11]}), .o(n441));   // memory_op.v(73)
    Mux_4u_16u Mux_441 (.sel({r1_op_inner}), .data({sys_r_addr[10], sys_r_addr[10], 
            sys_r_addr[10], sys_r_addr[10], sys_r_addr[10], r2[10], 
            a2[10], a1[10], sys_r_addr[10], sys_r_addr[10], sys_r_addr[10], 
            sys_r_addr[10], sys_r_addr[10], sys_r_addr[10], sys_r_addr[10], 
            sys_r_addr[10]}), .o(n442));   // memory_op.v(73)
    Mux_4u_16u Mux_442 (.sel({r1_op_inner}), .data({sys_r_addr[9], sys_r_addr[9], 
            sys_r_addr[9], sys_r_addr[9], sys_r_addr[9], r2[9], a2[9], 
            a1[9], sys_r_addr[9], sys_r_addr[9], sys_r_addr[9], sys_r_addr[9], 
            sys_r_addr[9], sys_r_addr[9], sys_r_addr[9], sys_r_addr[9]}), 
            .o(n443));   // memory_op.v(73)
    Mux_4u_16u Mux_443 (.sel({r1_op_inner}), .data({sys_r_addr[8], sys_r_addr[8], 
            sys_r_addr[8], sys_r_addr[8], sys_r_addr[8], r2[8], a2[8], 
            a1[8], sys_r_addr[8], sys_r_addr[8], sys_r_addr[8], sys_r_addr[8], 
            sys_r_addr[8], sys_r_addr[8], sys_r_addr[8], sys_r_addr[8]}), 
            .o(n444));   // memory_op.v(73)
    Mux_4u_16u Mux_444 (.sel({r1_op_inner}), .data({sys_r_addr[7], sys_r_addr[7], 
            sys_r_addr[7], sys_r_addr[7], sys_r_addr[7], r2[7], a2[7], 
            a1[7], sys_r_addr[7], sys_r_addr[7], sys_r_addr[7], sys_r_addr[7], 
            sys_r_addr[7], sys_r_addr[7], sys_r_addr[7], sys_r_addr[7]}), 
            .o(n445));   // memory_op.v(73)
    Mux_4u_16u Mux_445 (.sel({r1_op_inner}), .data({sys_r_addr[6], sys_r_addr[6], 
            sys_r_addr[6], sys_r_addr[6], sys_r_addr[6], r2[6], a2[6], 
            a1[6], sys_r_addr[6], sys_r_addr[6], sys_r_addr[6], sys_r_addr[6], 
            sys_r_addr[6], sys_r_addr[6], sys_r_addr[6], sys_r_addr[6]}), 
            .o(n446));   // memory_op.v(73)
    Mux_4u_16u Mux_446 (.sel({r1_op_inner}), .data({sys_r_addr[5], sys_r_addr[5], 
            sys_r_addr[5], sys_r_addr[5], sys_r_addr[5], r2[5], a2[5], 
            a1[5], sys_r_addr[5], sys_r_addr[5], sys_r_addr[5], sys_r_addr[5], 
            sys_r_addr[5], sys_r_addr[5], sys_r_addr[5], sys_r_addr[5]}), 
            .o(n447));   // memory_op.v(73)
    Mux_4u_16u Mux_447 (.sel({r1_op_inner}), .data({sys_r_addr[4], sys_r_addr[4], 
            sys_r_addr[4], sys_r_addr[4], sys_r_addr[4], r2[4], a2[4], 
            a1[4], sys_r_addr[4], sys_r_addr[4], sys_r_addr[4], sys_r_addr[4], 
            sys_r_addr[4], sys_r_addr[4], sys_r_addr[4], sys_r_addr[4]}), 
            .o(n448));   // memory_op.v(73)
    Mux_4u_16u Mux_448 (.sel({r1_op_inner}), .data({sys_r_addr[3], sys_r_addr[3], 
            sys_r_addr[3], sys_r_addr[3], sys_r_addr[3], r2[3], a2[3], 
            a1[3], sys_r_addr[3], sys_r_addr[3], sys_r_addr[3], sys_r_addr[3], 
            sys_r_addr[3], sys_r_addr[3], sys_r_addr[3], sys_r_addr[3]}), 
            .o(n449));   // memory_op.v(73)
    Mux_4u_16u Mux_449 (.sel({r1_op_inner}), .data({sys_r_addr[2], sys_r_addr[2], 
            sys_r_addr[2], sys_r_addr[2], sys_r_addr[2], r2[2], a2[2], 
            a1[2], sys_r_addr[2], sys_r_addr[2], sys_r_addr[2], sys_r_addr[2], 
            sys_r_addr[2], sys_r_addr[2], sys_r_addr[2], sys_r_addr[2]}), 
            .o(n450));   // memory_op.v(73)
    Mux_4u_16u Mux_450 (.sel({r1_op_inner}), .data({sys_r_addr[1], sys_r_addr[1], 
            sys_r_addr[1], sys_r_addr[1], sys_r_addr[1], r2[1], a2[1], 
            a1[1], sys_r_addr[1], sys_r_addr[1], sys_r_addr[1], sys_r_addr[1], 
            sys_r_addr[1], sys_r_addr[1], sys_r_addr[1], sys_r_addr[1]}), 
            .o(n451));   // memory_op.v(73)
    Mux_4u_16u Mux_451 (.sel({r1_op_inner}), .data({sys_r_addr[0], sys_r_addr[0], 
            sys_r_addr[0], sys_r_addr[0], sys_r_addr[0], r2[0], a2[0], 
            a1[0], sys_r_addr[0], sys_r_addr[0], sys_r_addr[0], sys_r_addr[0], 
            sys_r_addr[0], sys_r_addr[0], sys_r_addr[0], sys_r_addr[0]}), 
            .o(n452));   // memory_op.v(73)
    Mux_4u_16u Mux_452 (.sel({r1_op_inner}), .data({16'b0000011100000000}), 
            .o(n453));   // memory_op.v(73)
    Mux_4u_16u Mux_453 (.sel({r1_op_inner}), .data({ram_w_line[31], ram_w_line[31], 
            ram_w_line[31], ram_w_line[31], ram_w_line[31], ram_w_line[31], 
            ram_w_line[31], ram_w_line[31], r1[31], r1[31], r1[31], 
            ram_w_line[31], ram_w_line[31], ram_w_line[31], ram_w_line[31], 
            ram_w_line[31]}), .o(n454));   // memory_op.v(73)
    Mux_4u_16u Mux_454 (.sel({r1_op_inner}), .data({ram_w_line[30], ram_w_line[30], 
            ram_w_line[30], ram_w_line[30], ram_w_line[30], ram_w_line[30], 
            ram_w_line[30], ram_w_line[30], r1[30], r1[30], r1[30], 
            ram_w_line[30], ram_w_line[30], ram_w_line[30], ram_w_line[30], 
            ram_w_line[30]}), .o(n455));   // memory_op.v(73)
    Mux_4u_16u Mux_455 (.sel({r1_op_inner}), .data({ram_w_line[29], ram_w_line[29], 
            ram_w_line[29], ram_w_line[29], ram_w_line[29], ram_w_line[29], 
            ram_w_line[29], ram_w_line[29], r1[29], r1[29], r1[29], 
            ram_w_line[29], ram_w_line[29], ram_w_line[29], ram_w_line[29], 
            ram_w_line[29]}), .o(n456));   // memory_op.v(73)
    Mux_4u_16u Mux_456 (.sel({r1_op_inner}), .data({ram_w_line[28], ram_w_line[28], 
            ram_w_line[28], ram_w_line[28], ram_w_line[28], ram_w_line[28], 
            ram_w_line[28], ram_w_line[28], r1[28], r1[28], r1[28], 
            ram_w_line[28], ram_w_line[28], ram_w_line[28], ram_w_line[28], 
            ram_w_line[28]}), .o(n457));   // memory_op.v(73)
    Mux_4u_16u Mux_457 (.sel({r1_op_inner}), .data({ram_w_line[27], ram_w_line[27], 
            ram_w_line[27], ram_w_line[27], ram_w_line[27], ram_w_line[27], 
            ram_w_line[27], ram_w_line[27], r1[27], r1[27], r1[27], 
            ram_w_line[27], ram_w_line[27], ram_w_line[27], ram_w_line[27], 
            ram_w_line[27]}), .o(n458));   // memory_op.v(73)
    Mux_4u_16u Mux_458 (.sel({r1_op_inner}), .data({ram_w_line[26], ram_w_line[26], 
            ram_w_line[26], ram_w_line[26], ram_w_line[26], ram_w_line[26], 
            ram_w_line[26], ram_w_line[26], r1[26], r1[26], r1[26], 
            ram_w_line[26], ram_w_line[26], ram_w_line[26], ram_w_line[26], 
            ram_w_line[26]}), .o(n459));   // memory_op.v(73)
    Mux_4u_16u Mux_459 (.sel({r1_op_inner}), .data({ram_w_line[25], ram_w_line[25], 
            ram_w_line[25], ram_w_line[25], ram_w_line[25], ram_w_line[25], 
            ram_w_line[25], ram_w_line[25], r1[25], r1[25], r1[25], 
            ram_w_line[25], ram_w_line[25], ram_w_line[25], ram_w_line[25], 
            ram_w_line[25]}), .o(n460));   // memory_op.v(73)
    Mux_4u_16u Mux_460 (.sel({r1_op_inner}), .data({ram_w_line[24], ram_w_line[24], 
            ram_w_line[24], ram_w_line[24], ram_w_line[24], ram_w_line[24], 
            ram_w_line[24], ram_w_line[24], r1[24], r1[24], r1[24], 
            ram_w_line[24], ram_w_line[24], ram_w_line[24], ram_w_line[24], 
            ram_w_line[24]}), .o(n461));   // memory_op.v(73)
    Mux_4u_16u Mux_461 (.sel({r1_op_inner}), .data({ram_w_line[23], ram_w_line[23], 
            ram_w_line[23], ram_w_line[23], ram_w_line[23], ram_w_line[23], 
            ram_w_line[23], ram_w_line[23], r1[23], r1[23], r1[23], 
            ram_w_line[23], ram_w_line[23], ram_w_line[23], ram_w_line[23], 
            ram_w_line[23]}), .o(n462));   // memory_op.v(73)
    Mux_4u_16u Mux_462 (.sel({r1_op_inner}), .data({ram_w_line[22], ram_w_line[22], 
            ram_w_line[22], ram_w_line[22], ram_w_line[22], ram_w_line[22], 
            ram_w_line[22], ram_w_line[22], r1[22], r1[22], r1[22], 
            ram_w_line[22], ram_w_line[22], ram_w_line[22], ram_w_line[22], 
            ram_w_line[22]}), .o(n463));   // memory_op.v(73)
    Mux_4u_16u Mux_463 (.sel({r1_op_inner}), .data({ram_w_line[21], ram_w_line[21], 
            ram_w_line[21], ram_w_line[21], ram_w_line[21], ram_w_line[21], 
            ram_w_line[21], ram_w_line[21], r1[21], r1[21], r1[21], 
            ram_w_line[21], ram_w_line[21], ram_w_line[21], ram_w_line[21], 
            ram_w_line[21]}), .o(n464));   // memory_op.v(73)
    Mux_4u_16u Mux_464 (.sel({r1_op_inner}), .data({ram_w_line[20], ram_w_line[20], 
            ram_w_line[20], ram_w_line[20], ram_w_line[20], ram_w_line[20], 
            ram_w_line[20], ram_w_line[20], r1[20], r1[20], r1[20], 
            ram_w_line[20], ram_w_line[20], ram_w_line[20], ram_w_line[20], 
            ram_w_line[20]}), .o(n465));   // memory_op.v(73)
    Mux_4u_16u Mux_465 (.sel({r1_op_inner}), .data({ram_w_line[19], ram_w_line[19], 
            ram_w_line[19], ram_w_line[19], ram_w_line[19], ram_w_line[19], 
            ram_w_line[19], ram_w_line[19], r1[19], r1[19], r1[19], 
            ram_w_line[19], ram_w_line[19], ram_w_line[19], ram_w_line[19], 
            ram_w_line[19]}), .o(n466));   // memory_op.v(73)
    Mux_4u_16u Mux_466 (.sel({r1_op_inner}), .data({ram_w_line[18], ram_w_line[18], 
            ram_w_line[18], ram_w_line[18], ram_w_line[18], ram_w_line[18], 
            ram_w_line[18], ram_w_line[18], r1[18], r1[18], r1[18], 
            ram_w_line[18], ram_w_line[18], ram_w_line[18], ram_w_line[18], 
            ram_w_line[18]}), .o(n467));   // memory_op.v(73)
    Mux_4u_16u Mux_467 (.sel({r1_op_inner}), .data({ram_w_line[17], ram_w_line[17], 
            ram_w_line[17], ram_w_line[17], ram_w_line[17], ram_w_line[17], 
            ram_w_line[17], ram_w_line[17], r1[17], r1[17], r1[17], 
            ram_w_line[17], ram_w_line[17], ram_w_line[17], ram_w_line[17], 
            ram_w_line[17]}), .o(n468));   // memory_op.v(73)
    Mux_4u_16u Mux_468 (.sel({r1_op_inner}), .data({ram_w_line[16], ram_w_line[16], 
            ram_w_line[16], ram_w_line[16], ram_w_line[16], ram_w_line[16], 
            ram_w_line[16], ram_w_line[16], r1[16], r1[16], r1[16], 
            ram_w_line[16], ram_w_line[16], ram_w_line[16], ram_w_line[16], 
            ram_w_line[16]}), .o(n469));   // memory_op.v(73)
    Mux_4u_16u Mux_469 (.sel({r1_op_inner}), .data({ram_w_line[15], ram_w_line[15], 
            ram_w_line[15], ram_w_line[15], ram_w_line[15], ram_w_line[15], 
            ram_w_line[15], ram_w_line[15], r1[15], r1[15], r1[15], 
            ram_w_line[15], ram_w_line[15], ram_w_line[15], ram_w_line[15], 
            ram_w_line[15]}), .o(n470));   // memory_op.v(73)
    Mux_4u_16u Mux_470 (.sel({r1_op_inner}), .data({ram_w_line[14], ram_w_line[14], 
            ram_w_line[14], ram_w_line[14], ram_w_line[14], ram_w_line[14], 
            ram_w_line[14], ram_w_line[14], r1[14], r1[14], r1[14], 
            ram_w_line[14], ram_w_line[14], ram_w_line[14], ram_w_line[14], 
            ram_w_line[14]}), .o(n471));   // memory_op.v(73)
    Mux_4u_16u Mux_471 (.sel({r1_op_inner}), .data({ram_w_line[13], ram_w_line[13], 
            ram_w_line[13], ram_w_line[13], ram_w_line[13], ram_w_line[13], 
            ram_w_line[13], ram_w_line[13], r1[13], r1[13], r1[13], 
            ram_w_line[13], ram_w_line[13], ram_w_line[13], ram_w_line[13], 
            ram_w_line[13]}), .o(n472));   // memory_op.v(73)
    Mux_4u_16u Mux_472 (.sel({r1_op_inner}), .data({ram_w_line[12], ram_w_line[12], 
            ram_w_line[12], ram_w_line[12], ram_w_line[12], ram_w_line[12], 
            ram_w_line[12], ram_w_line[12], r1[12], r1[12], r1[12], 
            ram_w_line[12], ram_w_line[12], ram_w_line[12], ram_w_line[12], 
            ram_w_line[12]}), .o(n473));   // memory_op.v(73)
    Mux_4u_16u Mux_473 (.sel({r1_op_inner}), .data({ram_w_line[11], ram_w_line[11], 
            ram_w_line[11], ram_w_line[11], ram_w_line[11], ram_w_line[11], 
            ram_w_line[11], ram_w_line[11], r1[11], r1[11], r1[11], 
            ram_w_line[11], ram_w_line[11], ram_w_line[11], ram_w_line[11], 
            ram_w_line[11]}), .o(n474));   // memory_op.v(73)
    Mux_4u_16u Mux_474 (.sel({r1_op_inner}), .data({ram_w_line[10], ram_w_line[10], 
            ram_w_line[10], ram_w_line[10], ram_w_line[10], ram_w_line[10], 
            ram_w_line[10], ram_w_line[10], r1[10], r1[10], r1[10], 
            ram_w_line[10], ram_w_line[10], ram_w_line[10], ram_w_line[10], 
            ram_w_line[10]}), .o(n475));   // memory_op.v(73)
    Mux_4u_16u Mux_475 (.sel({r1_op_inner}), .data({ram_w_line[9], ram_w_line[9], 
            ram_w_line[9], ram_w_line[9], ram_w_line[9], ram_w_line[9], 
            ram_w_line[9], ram_w_line[9], r1[9], r1[9], r1[9], ram_w_line[9], 
            ram_w_line[9], ram_w_line[9], ram_w_line[9], ram_w_line[9]}), 
            .o(n476));   // memory_op.v(73)
    Mux_4u_16u Mux_476 (.sel({r1_op_inner}), .data({ram_w_line[8], ram_w_line[8], 
            ram_w_line[8], ram_w_line[8], ram_w_line[8], ram_w_line[8], 
            ram_w_line[8], ram_w_line[8], r1[8], r1[8], r1[8], ram_w_line[8], 
            ram_w_line[8], ram_w_line[8], ram_w_line[8], ram_w_line[8]}), 
            .o(n477));   // memory_op.v(73)
    Mux_4u_16u Mux_477 (.sel({r1_op_inner}), .data({ram_w_line[7], ram_w_line[7], 
            ram_w_line[7], ram_w_line[7], ram_w_line[7], ram_w_line[7], 
            ram_w_line[7], ram_w_line[7], r1[7], r1[7], r1[7], ram_w_line[7], 
            ram_w_line[7], ram_w_line[7], ram_w_line[7], ram_w_line[7]}), 
            .o(n478));   // memory_op.v(73)
    Mux_4u_16u Mux_478 (.sel({r1_op_inner}), .data({ram_w_line[6], ram_w_line[6], 
            ram_w_line[6], ram_w_line[6], ram_w_line[6], ram_w_line[6], 
            ram_w_line[6], ram_w_line[6], r1[6], r1[6], r1[6], ram_w_line[6], 
            ram_w_line[6], ram_w_line[6], ram_w_line[6], ram_w_line[6]}), 
            .o(n479));   // memory_op.v(73)
    Mux_4u_16u Mux_479 (.sel({r1_op_inner}), .data({ram_w_line[5], ram_w_line[5], 
            ram_w_line[5], ram_w_line[5], ram_w_line[5], ram_w_line[5], 
            ram_w_line[5], ram_w_line[5], r1[5], r1[5], r1[5], ram_w_line[5], 
            ram_w_line[5], ram_w_line[5], ram_w_line[5], ram_w_line[5]}), 
            .o(n480));   // memory_op.v(73)
    Mux_4u_16u Mux_480 (.sel({r1_op_inner}), .data({ram_w_line[4], ram_w_line[4], 
            ram_w_line[4], ram_w_line[4], ram_w_line[4], ram_w_line[4], 
            ram_w_line[4], ram_w_line[4], r1[4], r1[4], r1[4], ram_w_line[4], 
            ram_w_line[4], ram_w_line[4], ram_w_line[4], ram_w_line[4]}), 
            .o(n481));   // memory_op.v(73)
    Mux_4u_16u Mux_481 (.sel({r1_op_inner}), .data({ram_w_line[3], ram_w_line[3], 
            ram_w_line[3], ram_w_line[3], ram_w_line[3], ram_w_line[3], 
            ram_w_line[3], ram_w_line[3], r1[3], r1[3], r1[3], ram_w_line[3], 
            ram_w_line[3], ram_w_line[3], ram_w_line[3], ram_w_line[3]}), 
            .o(n482));   // memory_op.v(73)
    Mux_4u_16u Mux_482 (.sel({r1_op_inner}), .data({ram_w_line[2], ram_w_line[2], 
            ram_w_line[2], ram_w_line[2], ram_w_line[2], ram_w_line[2], 
            ram_w_line[2], ram_w_line[2], r1[2], r1[2], r1[2], ram_w_line[2], 
            ram_w_line[2], ram_w_line[2], ram_w_line[2], ram_w_line[2]}), 
            .o(n483));   // memory_op.v(73)
    Mux_4u_16u Mux_483 (.sel({r1_op_inner}), .data({ram_w_line[1], ram_w_line[1], 
            ram_w_line[1], ram_w_line[1], ram_w_line[1], ram_w_line[1], 
            ram_w_line[1], ram_w_line[1], r1[1], r1[1], r1[1], ram_w_line[1], 
            ram_w_line[1], ram_w_line[1], ram_w_line[1], ram_w_line[1]}), 
            .o(n484));   // memory_op.v(73)
    Mux_4u_16u Mux_484 (.sel({r1_op_inner}), .data({ram_w_line[0], ram_w_line[0], 
            ram_w_line[0], ram_w_line[0], ram_w_line[0], ram_w_line[0], 
            ram_w_line[0], ram_w_line[0], r1[0], r1[0], r1[0], ram_w_line[0], 
            ram_w_line[0], ram_w_line[0], ram_w_line[0], ram_w_line[0]}), 
            .o(n485));   // memory_op.v(73)
    Mux_4u_16u Mux_485 (.sel({r1_op_inner}), .data({ram_w_addr[31], ram_w_addr[31], 
            ram_w_addr[31], ram_w_addr[31], ram_w_addr[31], ram_w_addr[31], 
            ram_w_addr[31], ram_w_addr[31], r2[31], a2[31], a1[31], 
            ram_w_addr[31], ram_w_addr[31], ram_w_addr[31], ram_w_addr[31], 
            ram_w_addr[31]}), .o(n486));   // memory_op.v(73)
    Mux_4u_16u Mux_486 (.sel({r1_op_inner}), .data({ram_w_addr[30], ram_w_addr[30], 
            ram_w_addr[30], ram_w_addr[30], ram_w_addr[30], ram_w_addr[30], 
            ram_w_addr[30], ram_w_addr[30], r2[30], a2[30], a1[30], 
            ram_w_addr[30], ram_w_addr[30], ram_w_addr[30], ram_w_addr[30], 
            ram_w_addr[30]}), .o(n487));   // memory_op.v(73)
    Mux_4u_16u Mux_487 (.sel({r1_op_inner}), .data({ram_w_addr[29], ram_w_addr[29], 
            ram_w_addr[29], ram_w_addr[29], ram_w_addr[29], ram_w_addr[29], 
            ram_w_addr[29], ram_w_addr[29], r2[29], a2[29], a1[29], 
            ram_w_addr[29], ram_w_addr[29], ram_w_addr[29], ram_w_addr[29], 
            ram_w_addr[29]}), .o(n488));   // memory_op.v(73)
    Mux_4u_16u Mux_488 (.sel({r1_op_inner}), .data({ram_w_addr[28], ram_w_addr[28], 
            ram_w_addr[28], ram_w_addr[28], ram_w_addr[28], ram_w_addr[28], 
            ram_w_addr[28], ram_w_addr[28], r2[28], a2[28], a1[28], 
            ram_w_addr[28], ram_w_addr[28], ram_w_addr[28], ram_w_addr[28], 
            ram_w_addr[28]}), .o(n489));   // memory_op.v(73)
    Mux_4u_16u Mux_489 (.sel({r1_op_inner}), .data({ram_w_addr[27], ram_w_addr[27], 
            ram_w_addr[27], ram_w_addr[27], ram_w_addr[27], ram_w_addr[27], 
            ram_w_addr[27], ram_w_addr[27], r2[27], a2[27], a1[27], 
            ram_w_addr[27], ram_w_addr[27], ram_w_addr[27], ram_w_addr[27], 
            ram_w_addr[27]}), .o(n490));   // memory_op.v(73)
    Mux_4u_16u Mux_490 (.sel({r1_op_inner}), .data({ram_w_addr[26], ram_w_addr[26], 
            ram_w_addr[26], ram_w_addr[26], ram_w_addr[26], ram_w_addr[26], 
            ram_w_addr[26], ram_w_addr[26], r2[26], a2[26], a1[26], 
            ram_w_addr[26], ram_w_addr[26], ram_w_addr[26], ram_w_addr[26], 
            ram_w_addr[26]}), .o(n491));   // memory_op.v(73)
    Mux_4u_16u Mux_491 (.sel({r1_op_inner}), .data({ram_w_addr[25], ram_w_addr[25], 
            ram_w_addr[25], ram_w_addr[25], ram_w_addr[25], ram_w_addr[25], 
            ram_w_addr[25], ram_w_addr[25], r2[25], a2[25], a1[25], 
            ram_w_addr[25], ram_w_addr[25], ram_w_addr[25], ram_w_addr[25], 
            ram_w_addr[25]}), .o(n492));   // memory_op.v(73)
    Mux_4u_16u Mux_492 (.sel({r1_op_inner}), .data({ram_w_addr[24], ram_w_addr[24], 
            ram_w_addr[24], ram_w_addr[24], ram_w_addr[24], ram_w_addr[24], 
            ram_w_addr[24], ram_w_addr[24], r2[24], a2[24], a1[24], 
            ram_w_addr[24], ram_w_addr[24], ram_w_addr[24], ram_w_addr[24], 
            ram_w_addr[24]}), .o(n493));   // memory_op.v(73)
    Mux_4u_16u Mux_493 (.sel({r1_op_inner}), .data({ram_w_addr[23], ram_w_addr[23], 
            ram_w_addr[23], ram_w_addr[23], ram_w_addr[23], ram_w_addr[23], 
            ram_w_addr[23], ram_w_addr[23], r2[23], a2[23], a1[23], 
            ram_w_addr[23], ram_w_addr[23], ram_w_addr[23], ram_w_addr[23], 
            ram_w_addr[23]}), .o(n494));   // memory_op.v(73)
    Mux_4u_16u Mux_494 (.sel({r1_op_inner}), .data({ram_w_addr[22], ram_w_addr[22], 
            ram_w_addr[22], ram_w_addr[22], ram_w_addr[22], ram_w_addr[22], 
            ram_w_addr[22], ram_w_addr[22], r2[22], a2[22], a1[22], 
            ram_w_addr[22], ram_w_addr[22], ram_w_addr[22], ram_w_addr[22], 
            ram_w_addr[22]}), .o(n495));   // memory_op.v(73)
    Mux_4u_16u Mux_495 (.sel({r1_op_inner}), .data({ram_w_addr[21], ram_w_addr[21], 
            ram_w_addr[21], ram_w_addr[21], ram_w_addr[21], ram_w_addr[21], 
            ram_w_addr[21], ram_w_addr[21], r2[21], a2[21], a1[21], 
            ram_w_addr[21], ram_w_addr[21], ram_w_addr[21], ram_w_addr[21], 
            ram_w_addr[21]}), .o(n496));   // memory_op.v(73)
    Mux_4u_16u Mux_496 (.sel({r1_op_inner}), .data({ram_w_addr[20], ram_w_addr[20], 
            ram_w_addr[20], ram_w_addr[20], ram_w_addr[20], ram_w_addr[20], 
            ram_w_addr[20], ram_w_addr[20], r2[20], a2[20], a1[20], 
            ram_w_addr[20], ram_w_addr[20], ram_w_addr[20], ram_w_addr[20], 
            ram_w_addr[20]}), .o(n497));   // memory_op.v(73)
    Mux_4u_16u Mux_497 (.sel({r1_op_inner}), .data({ram_w_addr[19], ram_w_addr[19], 
            ram_w_addr[19], ram_w_addr[19], ram_w_addr[19], ram_w_addr[19], 
            ram_w_addr[19], ram_w_addr[19], r2[19], a2[19], a1[19], 
            ram_w_addr[19], ram_w_addr[19], ram_w_addr[19], ram_w_addr[19], 
            ram_w_addr[19]}), .o(n498));   // memory_op.v(73)
    Mux_4u_16u Mux_498 (.sel({r1_op_inner}), .data({ram_w_addr[18], ram_w_addr[18], 
            ram_w_addr[18], ram_w_addr[18], ram_w_addr[18], ram_w_addr[18], 
            ram_w_addr[18], ram_w_addr[18], r2[18], a2[18], a1[18], 
            ram_w_addr[18], ram_w_addr[18], ram_w_addr[18], ram_w_addr[18], 
            ram_w_addr[18]}), .o(n499));   // memory_op.v(73)
    Mux_4u_16u Mux_499 (.sel({r1_op_inner}), .data({ram_w_addr[17], ram_w_addr[17], 
            ram_w_addr[17], ram_w_addr[17], ram_w_addr[17], ram_w_addr[17], 
            ram_w_addr[17], ram_w_addr[17], r2[17], a2[17], a1[17], 
            ram_w_addr[17], ram_w_addr[17], ram_w_addr[17], ram_w_addr[17], 
            ram_w_addr[17]}), .o(n500));   // memory_op.v(73)
    Mux_4u_16u Mux_500 (.sel({r1_op_inner}), .data({ram_w_addr[16], ram_w_addr[16], 
            ram_w_addr[16], ram_w_addr[16], ram_w_addr[16], ram_w_addr[16], 
            ram_w_addr[16], ram_w_addr[16], r2[16], a2[16], a1[16], 
            ram_w_addr[16], ram_w_addr[16], ram_w_addr[16], ram_w_addr[16], 
            ram_w_addr[16]}), .o(n501));   // memory_op.v(73)
    Mux_4u_16u Mux_501 (.sel({r1_op_inner}), .data({ram_w_addr[15], ram_w_addr[15], 
            ram_w_addr[15], ram_w_addr[15], ram_w_addr[15], ram_w_addr[15], 
            ram_w_addr[15], ram_w_addr[15], r2[15], a2[15], a1[15], 
            ram_w_addr[15], ram_w_addr[15], ram_w_addr[15], ram_w_addr[15], 
            ram_w_addr[15]}), .o(n502));   // memory_op.v(73)
    Mux_4u_16u Mux_502 (.sel({r1_op_inner}), .data({ram_w_addr[14], ram_w_addr[14], 
            ram_w_addr[14], ram_w_addr[14], ram_w_addr[14], ram_w_addr[14], 
            ram_w_addr[14], ram_w_addr[14], r2[14], a2[14], a1[14], 
            ram_w_addr[14], ram_w_addr[14], ram_w_addr[14], ram_w_addr[14], 
            ram_w_addr[14]}), .o(n503));   // memory_op.v(73)
    Mux_4u_16u Mux_503 (.sel({r1_op_inner}), .data({ram_w_addr[13], ram_w_addr[13], 
            ram_w_addr[13], ram_w_addr[13], ram_w_addr[13], ram_w_addr[13], 
            ram_w_addr[13], ram_w_addr[13], r2[13], a2[13], a1[13], 
            ram_w_addr[13], ram_w_addr[13], ram_w_addr[13], ram_w_addr[13], 
            ram_w_addr[13]}), .o(n504));   // memory_op.v(73)
    Mux_4u_16u Mux_504 (.sel({r1_op_inner}), .data({ram_w_addr[12], ram_w_addr[12], 
            ram_w_addr[12], ram_w_addr[12], ram_w_addr[12], ram_w_addr[12], 
            ram_w_addr[12], ram_w_addr[12], r2[12], a2[12], a1[12], 
            ram_w_addr[12], ram_w_addr[12], ram_w_addr[12], ram_w_addr[12], 
            ram_w_addr[12]}), .o(n505));   // memory_op.v(73)
    Mux_4u_16u Mux_505 (.sel({r1_op_inner}), .data({ram_w_addr[11], ram_w_addr[11], 
            ram_w_addr[11], ram_w_addr[11], ram_w_addr[11], ram_w_addr[11], 
            ram_w_addr[11], ram_w_addr[11], r2[11], a2[11], a1[11], 
            ram_w_addr[11], ram_w_addr[11], ram_w_addr[11], ram_w_addr[11], 
            ram_w_addr[11]}), .o(n506));   // memory_op.v(73)
    Mux_4u_16u Mux_506 (.sel({r1_op_inner}), .data({ram_w_addr[10], ram_w_addr[10], 
            ram_w_addr[10], ram_w_addr[10], ram_w_addr[10], ram_w_addr[10], 
            ram_w_addr[10], ram_w_addr[10], r2[10], a2[10], a1[10], 
            ram_w_addr[10], ram_w_addr[10], ram_w_addr[10], ram_w_addr[10], 
            ram_w_addr[10]}), .o(n507));   // memory_op.v(73)
    Mux_4u_16u Mux_507 (.sel({r1_op_inner}), .data({ram_w_addr[9], ram_w_addr[9], 
            ram_w_addr[9], ram_w_addr[9], ram_w_addr[9], ram_w_addr[9], 
            ram_w_addr[9], ram_w_addr[9], r2[9], a2[9], a1[9], ram_w_addr[9], 
            ram_w_addr[9], ram_w_addr[9], ram_w_addr[9], ram_w_addr[9]}), 
            .o(n508));   // memory_op.v(73)
    Mux_4u_16u Mux_508 (.sel({r1_op_inner}), .data({ram_w_addr[8], ram_w_addr[8], 
            ram_w_addr[8], ram_w_addr[8], ram_w_addr[8], ram_w_addr[8], 
            ram_w_addr[8], ram_w_addr[8], r2[8], a2[8], a1[8], ram_w_addr[8], 
            ram_w_addr[8], ram_w_addr[8], ram_w_addr[8], ram_w_addr[8]}), 
            .o(n509));   // memory_op.v(73)
    Mux_4u_16u Mux_509 (.sel({r1_op_inner}), .data({ram_w_addr[7], ram_w_addr[7], 
            ram_w_addr[7], ram_w_addr[7], ram_w_addr[7], ram_w_addr[7], 
            ram_w_addr[7], ram_w_addr[7], r2[7], a2[7], a1[7], ram_w_addr[7], 
            ram_w_addr[7], ram_w_addr[7], ram_w_addr[7], ram_w_addr[7]}), 
            .o(n510));   // memory_op.v(73)
    Mux_4u_16u Mux_510 (.sel({r1_op_inner}), .data({ram_w_addr[6], ram_w_addr[6], 
            ram_w_addr[6], ram_w_addr[6], ram_w_addr[6], ram_w_addr[6], 
            ram_w_addr[6], ram_w_addr[6], r2[6], a2[6], a1[6], ram_w_addr[6], 
            ram_w_addr[6], ram_w_addr[6], ram_w_addr[6], ram_w_addr[6]}), 
            .o(n511));   // memory_op.v(73)
    Mux_4u_16u Mux_511 (.sel({r1_op_inner}), .data({ram_w_addr[5], ram_w_addr[5], 
            ram_w_addr[5], ram_w_addr[5], ram_w_addr[5], ram_w_addr[5], 
            ram_w_addr[5], ram_w_addr[5], r2[5], a2[5], a1[5], ram_w_addr[5], 
            ram_w_addr[5], ram_w_addr[5], ram_w_addr[5], ram_w_addr[5]}), 
            .o(n512));   // memory_op.v(73)
    Mux_4u_16u Mux_512 (.sel({r1_op_inner}), .data({ram_w_addr[4], ram_w_addr[4], 
            ram_w_addr[4], ram_w_addr[4], ram_w_addr[4], ram_w_addr[4], 
            ram_w_addr[4], ram_w_addr[4], r2[4], a2[4], a1[4], ram_w_addr[4], 
            ram_w_addr[4], ram_w_addr[4], ram_w_addr[4], ram_w_addr[4]}), 
            .o(n513));   // memory_op.v(73)
    Mux_4u_16u Mux_513 (.sel({r1_op_inner}), .data({ram_w_addr[3], ram_w_addr[3], 
            ram_w_addr[3], ram_w_addr[3], ram_w_addr[3], ram_w_addr[3], 
            ram_w_addr[3], ram_w_addr[3], r2[3], a2[3], a1[3], ram_w_addr[3], 
            ram_w_addr[3], ram_w_addr[3], ram_w_addr[3], ram_w_addr[3]}), 
            .o(n514));   // memory_op.v(73)
    Mux_4u_16u Mux_514 (.sel({r1_op_inner}), .data({ram_w_addr[2], ram_w_addr[2], 
            ram_w_addr[2], ram_w_addr[2], ram_w_addr[2], ram_w_addr[2], 
            ram_w_addr[2], ram_w_addr[2], r2[2], a2[2], a1[2], ram_w_addr[2], 
            ram_w_addr[2], ram_w_addr[2], ram_w_addr[2], ram_w_addr[2]}), 
            .o(n515));   // memory_op.v(73)
    Mux_4u_16u Mux_515 (.sel({r1_op_inner}), .data({ram_w_addr[1], ram_w_addr[1], 
            ram_w_addr[1], ram_w_addr[1], ram_w_addr[1], ram_w_addr[1], 
            ram_w_addr[1], ram_w_addr[1], r2[1], a2[1], a1[1], ram_w_addr[1], 
            ram_w_addr[1], ram_w_addr[1], ram_w_addr[1], ram_w_addr[1]}), 
            .o(n516));   // memory_op.v(73)
    Mux_4u_16u Mux_516 (.sel({r1_op_inner}), .data({ram_w_addr[0], ram_w_addr[0], 
            ram_w_addr[0], ram_w_addr[0], ram_w_addr[0], ram_w_addr[0], 
            ram_w_addr[0], ram_w_addr[0], r2[0], a2[0], a1[0], ram_w_addr[0], 
            ram_w_addr[0], ram_w_addr[0], ram_w_addr[0], ram_w_addr[0]}), 
            .o(n517));   // memory_op.v(73)
    Mux_4u_16u Mux_517 (.sel({r1_op_inner}), .data({16'b0000000011100000}), 
            .o(n518));   // memory_op.v(73)
    Mux_4u_16u Mux_518 (.sel({r1_op_inner}), .data({ram_r_addr[31], ram_r_addr[31], 
            ram_r_addr[31], ram_r_addr[31], ram_r_addr[31], ram_r_addr[31], 
            ram_r_addr[31], ram_r_addr[31], ram_r_addr[31], ram_r_addr[31], 
            ram_r_addr[31], r2[31], a2[31], a1[31], ram_r_addr[31], 
            ram_r_addr[31]}), .o(n519));   // memory_op.v(73)
    Mux_4u_16u Mux_519 (.sel({r1_op_inner}), .data({ram_r_addr[30], ram_r_addr[30], 
            ram_r_addr[30], ram_r_addr[30], ram_r_addr[30], ram_r_addr[30], 
            ram_r_addr[30], ram_r_addr[30], ram_r_addr[30], ram_r_addr[30], 
            ram_r_addr[30], r2[30], a2[30], a1[30], ram_r_addr[30], 
            ram_r_addr[30]}), .o(n520));   // memory_op.v(73)
    Mux_4u_16u Mux_520 (.sel({r1_op_inner}), .data({ram_r_addr[29], ram_r_addr[29], 
            ram_r_addr[29], ram_r_addr[29], ram_r_addr[29], ram_r_addr[29], 
            ram_r_addr[29], ram_r_addr[29], ram_r_addr[29], ram_r_addr[29], 
            ram_r_addr[29], r2[29], a2[29], a1[29], ram_r_addr[29], 
            ram_r_addr[29]}), .o(n521));   // memory_op.v(73)
    Mux_4u_16u Mux_521 (.sel({r1_op_inner}), .data({ram_r_addr[28], ram_r_addr[28], 
            ram_r_addr[28], ram_r_addr[28], ram_r_addr[28], ram_r_addr[28], 
            ram_r_addr[28], ram_r_addr[28], ram_r_addr[28], ram_r_addr[28], 
            ram_r_addr[28], r2[28], a2[28], a1[28], ram_r_addr[28], 
            ram_r_addr[28]}), .o(n522));   // memory_op.v(73)
    Mux_4u_16u Mux_522 (.sel({r1_op_inner}), .data({ram_r_addr[27], ram_r_addr[27], 
            ram_r_addr[27], ram_r_addr[27], ram_r_addr[27], ram_r_addr[27], 
            ram_r_addr[27], ram_r_addr[27], ram_r_addr[27], ram_r_addr[27], 
            ram_r_addr[27], r2[27], a2[27], a1[27], ram_r_addr[27], 
            ram_r_addr[27]}), .o(n523));   // memory_op.v(73)
    Mux_4u_16u Mux_523 (.sel({r1_op_inner}), .data({ram_r_addr[26], ram_r_addr[26], 
            ram_r_addr[26], ram_r_addr[26], ram_r_addr[26], ram_r_addr[26], 
            ram_r_addr[26], ram_r_addr[26], ram_r_addr[26], ram_r_addr[26], 
            ram_r_addr[26], r2[26], a2[26], a1[26], ram_r_addr[26], 
            ram_r_addr[26]}), .o(n524));   // memory_op.v(73)
    Mux_4u_16u Mux_524 (.sel({r1_op_inner}), .data({ram_r_addr[25], ram_r_addr[25], 
            ram_r_addr[25], ram_r_addr[25], ram_r_addr[25], ram_r_addr[25], 
            ram_r_addr[25], ram_r_addr[25], ram_r_addr[25], ram_r_addr[25], 
            ram_r_addr[25], r2[25], a2[25], a1[25], ram_r_addr[25], 
            ram_r_addr[25]}), .o(n525));   // memory_op.v(73)
    Mux_4u_16u Mux_525 (.sel({r1_op_inner}), .data({ram_r_addr[24], ram_r_addr[24], 
            ram_r_addr[24], ram_r_addr[24], ram_r_addr[24], ram_r_addr[24], 
            ram_r_addr[24], ram_r_addr[24], ram_r_addr[24], ram_r_addr[24], 
            ram_r_addr[24], r2[24], a2[24], a1[24], ram_r_addr[24], 
            ram_r_addr[24]}), .o(n526));   // memory_op.v(73)
    Mux_4u_16u Mux_526 (.sel({r1_op_inner}), .data({ram_r_addr[23], ram_r_addr[23], 
            ram_r_addr[23], ram_r_addr[23], ram_r_addr[23], ram_r_addr[23], 
            ram_r_addr[23], ram_r_addr[23], ram_r_addr[23], ram_r_addr[23], 
            ram_r_addr[23], r2[23], a2[23], a1[23], ram_r_addr[23], 
            ram_r_addr[23]}), .o(n527));   // memory_op.v(73)
    Mux_4u_16u Mux_527 (.sel({r1_op_inner}), .data({ram_r_addr[22], ram_r_addr[22], 
            ram_r_addr[22], ram_r_addr[22], ram_r_addr[22], ram_r_addr[22], 
            ram_r_addr[22], ram_r_addr[22], ram_r_addr[22], ram_r_addr[22], 
            ram_r_addr[22], r2[22], a2[22], a1[22], ram_r_addr[22], 
            ram_r_addr[22]}), .o(n528));   // memory_op.v(73)
    Mux_4u_16u Mux_528 (.sel({r1_op_inner}), .data({ram_r_addr[21], ram_r_addr[21], 
            ram_r_addr[21], ram_r_addr[21], ram_r_addr[21], ram_r_addr[21], 
            ram_r_addr[21], ram_r_addr[21], ram_r_addr[21], ram_r_addr[21], 
            ram_r_addr[21], r2[21], a2[21], a1[21], ram_r_addr[21], 
            ram_r_addr[21]}), .o(n529));   // memory_op.v(73)
    Mux_4u_16u Mux_529 (.sel({r1_op_inner}), .data({ram_r_addr[20], ram_r_addr[20], 
            ram_r_addr[20], ram_r_addr[20], ram_r_addr[20], ram_r_addr[20], 
            ram_r_addr[20], ram_r_addr[20], ram_r_addr[20], ram_r_addr[20], 
            ram_r_addr[20], r2[20], a2[20], a1[20], ram_r_addr[20], 
            ram_r_addr[20]}), .o(n530));   // memory_op.v(73)
    Mux_4u_16u Mux_530 (.sel({r1_op_inner}), .data({ram_r_addr[19], ram_r_addr[19], 
            ram_r_addr[19], ram_r_addr[19], ram_r_addr[19], ram_r_addr[19], 
            ram_r_addr[19], ram_r_addr[19], ram_r_addr[19], ram_r_addr[19], 
            ram_r_addr[19], r2[19], a2[19], a1[19], ram_r_addr[19], 
            ram_r_addr[19]}), .o(n531));   // memory_op.v(73)
    Mux_4u_16u Mux_531 (.sel({r1_op_inner}), .data({ram_r_addr[18], ram_r_addr[18], 
            ram_r_addr[18], ram_r_addr[18], ram_r_addr[18], ram_r_addr[18], 
            ram_r_addr[18], ram_r_addr[18], ram_r_addr[18], ram_r_addr[18], 
            ram_r_addr[18], r2[18], a2[18], a1[18], ram_r_addr[18], 
            ram_r_addr[18]}), .o(n532));   // memory_op.v(73)
    Mux_4u_16u Mux_532 (.sel({r1_op_inner}), .data({ram_r_addr[17], ram_r_addr[17], 
            ram_r_addr[17], ram_r_addr[17], ram_r_addr[17], ram_r_addr[17], 
            ram_r_addr[17], ram_r_addr[17], ram_r_addr[17], ram_r_addr[17], 
            ram_r_addr[17], r2[17], a2[17], a1[17], ram_r_addr[17], 
            ram_r_addr[17]}), .o(n533));   // memory_op.v(73)
    Mux_4u_16u Mux_533 (.sel({r1_op_inner}), .data({ram_r_addr[16], ram_r_addr[16], 
            ram_r_addr[16], ram_r_addr[16], ram_r_addr[16], ram_r_addr[16], 
            ram_r_addr[16], ram_r_addr[16], ram_r_addr[16], ram_r_addr[16], 
            ram_r_addr[16], r2[16], a2[16], a1[16], ram_r_addr[16], 
            ram_r_addr[16]}), .o(n534));   // memory_op.v(73)
    Mux_4u_16u Mux_534 (.sel({r1_op_inner}), .data({ram_r_addr[15], ram_r_addr[15], 
            ram_r_addr[15], ram_r_addr[15], ram_r_addr[15], ram_r_addr[15], 
            ram_r_addr[15], ram_r_addr[15], ram_r_addr[15], ram_r_addr[15], 
            ram_r_addr[15], r2[15], a2[15], a1[15], ram_r_addr[15], 
            ram_r_addr[15]}), .o(n535));   // memory_op.v(73)
    Mux_4u_16u Mux_535 (.sel({r1_op_inner}), .data({ram_r_addr[14], ram_r_addr[14], 
            ram_r_addr[14], ram_r_addr[14], ram_r_addr[14], ram_r_addr[14], 
            ram_r_addr[14], ram_r_addr[14], ram_r_addr[14], ram_r_addr[14], 
            ram_r_addr[14], r2[14], a2[14], a1[14], ram_r_addr[14], 
            ram_r_addr[14]}), .o(n536));   // memory_op.v(73)
    Mux_4u_16u Mux_536 (.sel({r1_op_inner}), .data({ram_r_addr[13], ram_r_addr[13], 
            ram_r_addr[13], ram_r_addr[13], ram_r_addr[13], ram_r_addr[13], 
            ram_r_addr[13], ram_r_addr[13], ram_r_addr[13], ram_r_addr[13], 
            ram_r_addr[13], r2[13], a2[13], a1[13], ram_r_addr[13], 
            ram_r_addr[13]}), .o(n537));   // memory_op.v(73)
    Mux_4u_16u Mux_537 (.sel({r1_op_inner}), .data({ram_r_addr[12], ram_r_addr[12], 
            ram_r_addr[12], ram_r_addr[12], ram_r_addr[12], ram_r_addr[12], 
            ram_r_addr[12], ram_r_addr[12], ram_r_addr[12], ram_r_addr[12], 
            ram_r_addr[12], r2[12], a2[12], a1[12], ram_r_addr[12], 
            ram_r_addr[12]}), .o(n538));   // memory_op.v(73)
    Mux_4u_16u Mux_538 (.sel({r1_op_inner}), .data({ram_r_addr[11], ram_r_addr[11], 
            ram_r_addr[11], ram_r_addr[11], ram_r_addr[11], ram_r_addr[11], 
            ram_r_addr[11], ram_r_addr[11], ram_r_addr[11], ram_r_addr[11], 
            ram_r_addr[11], r2[11], a2[11], a1[11], ram_r_addr[11], 
            ram_r_addr[11]}), .o(n539));   // memory_op.v(73)
    Mux_4u_16u Mux_539 (.sel({r1_op_inner}), .data({ram_r_addr[10], ram_r_addr[10], 
            ram_r_addr[10], ram_r_addr[10], ram_r_addr[10], ram_r_addr[10], 
            ram_r_addr[10], ram_r_addr[10], ram_r_addr[10], ram_r_addr[10], 
            ram_r_addr[10], r2[10], a2[10], a1[10], ram_r_addr[10], 
            ram_r_addr[10]}), .o(n540));   // memory_op.v(73)
    Mux_4u_16u Mux_540 (.sel({r1_op_inner}), .data({ram_r_addr[9], ram_r_addr[9], 
            ram_r_addr[9], ram_r_addr[9], ram_r_addr[9], ram_r_addr[9], 
            ram_r_addr[9], ram_r_addr[9], ram_r_addr[9], ram_r_addr[9], 
            ram_r_addr[9], r2[9], a2[9], a1[9], ram_r_addr[9], ram_r_addr[9]}), 
            .o(n541));   // memory_op.v(73)
    Mux_4u_16u Mux_541 (.sel({r1_op_inner}), .data({ram_r_addr[8], ram_r_addr[8], 
            ram_r_addr[8], ram_r_addr[8], ram_r_addr[8], ram_r_addr[8], 
            ram_r_addr[8], ram_r_addr[8], ram_r_addr[8], ram_r_addr[8], 
            ram_r_addr[8], r2[8], a2[8], a1[8], ram_r_addr[8], ram_r_addr[8]}), 
            .o(n542));   // memory_op.v(73)
    Mux_4u_16u Mux_542 (.sel({r1_op_inner}), .data({ram_r_addr[7], ram_r_addr[7], 
            ram_r_addr[7], ram_r_addr[7], ram_r_addr[7], ram_r_addr[7], 
            ram_r_addr[7], ram_r_addr[7], ram_r_addr[7], ram_r_addr[7], 
            ram_r_addr[7], r2[7], a2[7], a1[7], ram_r_addr[7], ram_r_addr[7]}), 
            .o(n543));   // memory_op.v(73)
    Mux_4u_16u Mux_543 (.sel({r1_op_inner}), .data({ram_r_addr[6], ram_r_addr[6], 
            ram_r_addr[6], ram_r_addr[6], ram_r_addr[6], ram_r_addr[6], 
            ram_r_addr[6], ram_r_addr[6], ram_r_addr[6], ram_r_addr[6], 
            ram_r_addr[6], r2[6], a2[6], a1[6], ram_r_addr[6], ram_r_addr[6]}), 
            .o(n544));   // memory_op.v(73)
    Mux_4u_16u Mux_544 (.sel({r1_op_inner}), .data({ram_r_addr[5], ram_r_addr[5], 
            ram_r_addr[5], ram_r_addr[5], ram_r_addr[5], ram_r_addr[5], 
            ram_r_addr[5], ram_r_addr[5], ram_r_addr[5], ram_r_addr[5], 
            ram_r_addr[5], r2[5], a2[5], a1[5], ram_r_addr[5], ram_r_addr[5]}), 
            .o(n545));   // memory_op.v(73)
    Mux_4u_16u Mux_545 (.sel({r1_op_inner}), .data({ram_r_addr[4], ram_r_addr[4], 
            ram_r_addr[4], ram_r_addr[4], ram_r_addr[4], ram_r_addr[4], 
            ram_r_addr[4], ram_r_addr[4], ram_r_addr[4], ram_r_addr[4], 
            ram_r_addr[4], r2[4], a2[4], a1[4], ram_r_addr[4], ram_r_addr[4]}), 
            .o(n546));   // memory_op.v(73)
    Mux_4u_16u Mux_546 (.sel({r1_op_inner}), .data({ram_r_addr[3], ram_r_addr[3], 
            ram_r_addr[3], ram_r_addr[3], ram_r_addr[3], ram_r_addr[3], 
            ram_r_addr[3], ram_r_addr[3], ram_r_addr[3], ram_r_addr[3], 
            ram_r_addr[3], r2[3], a2[3], a1[3], ram_r_addr[3], ram_r_addr[3]}), 
            .o(n547));   // memory_op.v(73)
    Mux_4u_16u Mux_547 (.sel({r1_op_inner}), .data({ram_r_addr[2], ram_r_addr[2], 
            ram_r_addr[2], ram_r_addr[2], ram_r_addr[2], ram_r_addr[2], 
            ram_r_addr[2], ram_r_addr[2], ram_r_addr[2], ram_r_addr[2], 
            ram_r_addr[2], r2[2], a2[2], a1[2], ram_r_addr[2], ram_r_addr[2]}), 
            .o(n548));   // memory_op.v(73)
    Mux_4u_16u Mux_548 (.sel({r1_op_inner}), .data({ram_r_addr[1], ram_r_addr[1], 
            ram_r_addr[1], ram_r_addr[1], ram_r_addr[1], ram_r_addr[1], 
            ram_r_addr[1], ram_r_addr[1], ram_r_addr[1], ram_r_addr[1], 
            ram_r_addr[1], r2[1], a2[1], a1[1], ram_r_addr[1], ram_r_addr[1]}), 
            .o(n549));   // memory_op.v(73)
    Mux_4u_16u Mux_549 (.sel({r1_op_inner}), .data({ram_r_addr[0], ram_r_addr[0], 
            ram_r_addr[0], ram_r_addr[0], ram_r_addr[0], ram_r_addr[0], 
            ram_r_addr[0], ram_r_addr[0], ram_r_addr[0], ram_r_addr[0], 
            ram_r_addr[0], r2[0], a2[0], a1[0], ram_r_addr[0], ram_r_addr[0]}), 
            .o(n550));   // memory_op.v(73)
    Mux_4u_16u Mux_550 (.sel({r1_op_inner}), .data({16'b0000000000011100}), 
            .o(n551));   // memory_op.v(73)
    Mux_4u_16u Mux_551 (.sel({r2_op_inner}), .data({m2_select[2], 15'b000011100000000}), 
            .o(n552));   // memory_op.v(166)
    Mux_4u_16u Mux_552 (.sel({r2_op_inner}), .data({m2_select[1], 15'b011100011111110}), 
            .o(n553));   // memory_op.v(166)
    Mux_4u_16u Mux_553 (.sel({r2_op_inner}), .data({m2_select[0], 15'b100000000011100}), 
            .o(n554));   // memory_op.v(166)
    Mux_4u_16u Mux_554 (.sel({r2_op_inner}), .data({n356, n356, r2[31], 
            r2[31], r2[31], n356, n356, n356, n356, n356, n356, 
            n356, n356, n356, n356, n356}), .o(n555));   // memory_op.v(166)
    Mux_4u_16u Mux_555 (.sel({r2_op_inner}), .data({n357, n357, r2[30], 
            r2[30], r2[30], n357, n357, n357, n357, n357, n357, 
            n357, n357, n357, n357, n357}), .o(n556));   // memory_op.v(166)
    Mux_4u_16u Mux_556 (.sel({r2_op_inner}), .data({n358, n358, r2[29], 
            r2[29], r2[29], n358, n358, n358, n358, n358, n358, 
            n358, n358, n358, n358, n358}), .o(n557));   // memory_op.v(166)
    Mux_4u_16u Mux_557 (.sel({r2_op_inner}), .data({n359, n359, r2[28], 
            r2[28], r2[28], n359, n359, n359, n359, n359, n359, 
            n359, n359, n359, n359, n359}), .o(n558));   // memory_op.v(166)
    Mux_4u_16u Mux_558 (.sel({r2_op_inner}), .data({n360, n360, r2[27], 
            r2[27], r2[27], n360, n360, n360, n360, n360, n360, 
            n360, n360, n360, n360, n360}), .o(n559));   // memory_op.v(166)
    Mux_4u_16u Mux_559 (.sel({r2_op_inner}), .data({n361, n361, r2[26], 
            r2[26], r2[26], n361, n361, n361, n361, n361, n361, 
            n361, n361, n361, n361, n361}), .o(n560));   // memory_op.v(166)
    Mux_4u_16u Mux_560 (.sel({r2_op_inner}), .data({n362, n362, r2[25], 
            r2[25], r2[25], n362, n362, n362, n362, n362, n362, 
            n362, n362, n362, n362, n362}), .o(n561));   // memory_op.v(166)
    Mux_4u_16u Mux_561 (.sel({r2_op_inner}), .data({n363, n363, r2[24], 
            r2[24], r2[24], n363, n363, n363, n363, n363, n363, 
            n363, n363, n363, n363, n363}), .o(n562));   // memory_op.v(166)
    Mux_4u_16u Mux_562 (.sel({r2_op_inner}), .data({n364, n364, r2[23], 
            r2[23], r2[23], n364, n364, n364, n364, n364, n364, 
            n364, n364, n364, n364, n364}), .o(n563));   // memory_op.v(166)
    Mux_4u_16u Mux_563 (.sel({r2_op_inner}), .data({n365, n365, r2[22], 
            r2[22], r2[22], n365, n365, n365, n365, n365, n365, 
            n365, n365, n365, n365, n365}), .o(n564));   // memory_op.v(166)
    Mux_4u_16u Mux_564 (.sel({r2_op_inner}), .data({n366, n366, r2[21], 
            r2[21], r2[21], n366, n366, n366, n366, n366, n366, 
            n366, n366, n366, n366, n366}), .o(n565));   // memory_op.v(166)
    Mux_4u_16u Mux_565 (.sel({r2_op_inner}), .data({n367, n367, r2[20], 
            r2[20], r2[20], n367, n367, n367, n367, n367, n367, 
            n367, n367, n367, n367, n367}), .o(n566));   // memory_op.v(166)
    Mux_4u_16u Mux_566 (.sel({r2_op_inner}), .data({n368, n368, r2[19], 
            r2[19], r2[19], n368, n368, n368, n368, n368, n368, 
            n368, n368, n368, n368, n368}), .o(n567));   // memory_op.v(166)
    Mux_4u_16u Mux_567 (.sel({r2_op_inner}), .data({n369, n369, r2[18], 
            r2[18], r2[18], n369, n369, n369, n369, n369, n369, 
            n369, n369, n369, n369, n369}), .o(n568));   // memory_op.v(166)
    Mux_4u_16u Mux_568 (.sel({r2_op_inner}), .data({n370, n370, r2[17], 
            r2[17], r2[17], n370, n370, n370, n370, n370, n370, 
            n370, n370, n370, n370, n370}), .o(n569));   // memory_op.v(166)
    Mux_4u_16u Mux_569 (.sel({r2_op_inner}), .data({n371, n371, r2[16], 
            r2[16], r2[16], n371, n371, n371, n371, n371, n371, 
            n371, n371, n371, n371, n371}), .o(n570));   // memory_op.v(166)
    Mux_4u_16u Mux_570 (.sel({r2_op_inner}), .data({n372, n372, r2[15], 
            r2[15], r2[15], n372, n372, n372, n372, n372, n372, 
            n372, n372, n372, n372, n372}), .o(n571));   // memory_op.v(166)
    Mux_4u_16u Mux_571 (.sel({r2_op_inner}), .data({n373, n373, r2[14], 
            r2[14], r2[14], n373, n373, n373, n373, n373, n373, 
            n373, n373, n373, n373, n373}), .o(n572));   // memory_op.v(166)
    Mux_4u_16u Mux_572 (.sel({r2_op_inner}), .data({n374, n374, r2[13], 
            r2[13], r2[13], n374, n374, n374, n374, n374, n374, 
            n374, n374, n374, n374, n374}), .o(n573));   // memory_op.v(166)
    Mux_4u_16u Mux_573 (.sel({r2_op_inner}), .data({n375, n375, r2[12], 
            r2[12], r2[12], n375, n375, n375, n375, n375, n375, 
            n375, n375, n375, n375, n375}), .o(n574));   // memory_op.v(166)
    Mux_4u_16u Mux_574 (.sel({r2_op_inner}), .data({n376, n376, r2[11], 
            r2[11], r2[11], n376, n376, n376, n376, n376, n376, 
            n376, n376, n376, n376, n376}), .o(n575));   // memory_op.v(166)
    Mux_4u_16u Mux_575 (.sel({r2_op_inner}), .data({n377, n377, r2[10], 
            r2[10], r2[10], n377, n377, n377, n377, n377, n377, 
            n377, n377, n377, n377, n377}), .o(n576));   // memory_op.v(166)
    Mux_4u_16u Mux_576 (.sel({r2_op_inner}), .data({n378, n378, r2[9], 
            r2[9], r2[9], n378, n378, n378, n378, n378, n378, 
            n378, n378, n378, n378, n378}), .o(n577));   // memory_op.v(166)
    Mux_4u_16u Mux_577 (.sel({r2_op_inner}), .data({n379, n379, r2[8], 
            r2[8], r2[8], n379, n379, n379, n379, n379, n379, 
            n379, n379, n379, n379, n379}), .o(n578));   // memory_op.v(166)
    Mux_4u_16u Mux_578 (.sel({r2_op_inner}), .data({n380, n380, r2[7], 
            r2[7], r2[7], n380, n380, n380, n380, n380, n380, 
            n380, n380, n380, n380, n380}), .o(n579));   // memory_op.v(166)
    Mux_4u_16u Mux_579 (.sel({r2_op_inner}), .data({n381, n381, r2[6], 
            r2[6], r2[6], n381, n381, n381, n381, n381, n381, 
            n381, n381, n381, n381, n381}), .o(n580));   // memory_op.v(166)
    Mux_4u_16u Mux_580 (.sel({r2_op_inner}), .data({n382, n382, r2[5], 
            r2[5], r2[5], n382, n382, n382, n382, n382, n382, 
            n382, n382, n382, n382, n382}), .o(n581));   // memory_op.v(166)
    Mux_4u_16u Mux_581 (.sel({r2_op_inner}), .data({n383, n383, r2[4], 
            r2[4], r2[4], n383, n383, n383, n383, n383, n383, 
            n383, n383, n383, n383, n383}), .o(n582));   // memory_op.v(166)
    Mux_4u_16u Mux_582 (.sel({r2_op_inner}), .data({n384, n384, r2[3], 
            r2[3], r2[3], n384, n384, n384, n384, n384, n384, 
            n384, n384, n384, n384, n384}), .o(n583));   // memory_op.v(166)
    Mux_4u_16u Mux_583 (.sel({r2_op_inner}), .data({n385, n385, r2[2], 
            r2[2], r2[2], n385, n385, n385, n385, n385, n385, 
            n385, n385, n385, n385, n385}), .o(n584));   // memory_op.v(166)
    Mux_4u_16u Mux_584 (.sel({r2_op_inner}), .data({n386, n386, r2[1], 
            r2[1], r2[1], n386, n386, n386, n386, n386, n386, 
            n386, n386, n386, n386, n386}), .o(n585));   // memory_op.v(166)
    Mux_4u_16u Mux_585 (.sel({r2_op_inner}), .data({n387, n387, r2[0], 
            r2[0], r2[0], n387, n387, n387, n387, n387, n387, 
            n387, n387, n387, n387, n387}), .o(n586));   // memory_op.v(166)
    Mux_4u_16u Mux_586 (.sel({r2_op_inner}), .data({n388, n388, r1[31], 
            a2[31], a1[31], n388, n388, n388, n388, n388, n388, 
            n388, n388, n388, n388, n388}), .o(n587));   // memory_op.v(166)
    Mux_4u_16u Mux_587 (.sel({r2_op_inner}), .data({n389, n389, r1[30], 
            a2[30], a1[30], n389, n389, n389, n389, n389, n389, 
            n389, n389, n389, n389, n389}), .o(n588));   // memory_op.v(166)
    Mux_4u_16u Mux_588 (.sel({r2_op_inner}), .data({n390, n390, r1[29], 
            a2[29], a1[29], n390, n390, n390, n390, n390, n390, 
            n390, n390, n390, n390, n390}), .o(n589));   // memory_op.v(166)
    Mux_4u_16u Mux_589 (.sel({r2_op_inner}), .data({n391, n391, r1[28], 
            a2[28], a1[28], n391, n391, n391, n391, n391, n391, 
            n391, n391, n391, n391, n391}), .o(n590));   // memory_op.v(166)
    Mux_4u_16u Mux_590 (.sel({r2_op_inner}), .data({n392, n392, r1[27], 
            a2[27], a1[27], n392, n392, n392, n392, n392, n392, 
            n392, n392, n392, n392, n392}), .o(n591));   // memory_op.v(166)
    Mux_4u_16u Mux_591 (.sel({r2_op_inner}), .data({n393, n393, r1[26], 
            a2[26], a1[26], n393, n393, n393, n393, n393, n393, 
            n393, n393, n393, n393, n393}), .o(n592));   // memory_op.v(166)
    Mux_4u_16u Mux_592 (.sel({r2_op_inner}), .data({n394, n394, r1[25], 
            a2[25], a1[25], n394, n394, n394, n394, n394, n394, 
            n394, n394, n394, n394, n394}), .o(n593));   // memory_op.v(166)
    Mux_4u_16u Mux_593 (.sel({r2_op_inner}), .data({n395, n395, r1[24], 
            a2[24], a1[24], n395, n395, n395, n395, n395, n395, 
            n395, n395, n395, n395, n395}), .o(n594));   // memory_op.v(166)
    Mux_4u_16u Mux_594 (.sel({r2_op_inner}), .data({n396, n396, r1[23], 
            a2[23], a1[23], n396, n396, n396, n396, n396, n396, 
            n396, n396, n396, n396, n396}), .o(n595));   // memory_op.v(166)
    Mux_4u_16u Mux_595 (.sel({r2_op_inner}), .data({n397, n397, r1[22], 
            a2[22], a1[22], n397, n397, n397, n397, n397, n397, 
            n397, n397, n397, n397, n397}), .o(n596));   // memory_op.v(166)
    Mux_4u_16u Mux_596 (.sel({r2_op_inner}), .data({n398, n398, r1[21], 
            a2[21], a1[21], n398, n398, n398, n398, n398, n398, 
            n398, n398, n398, n398, n398}), .o(n597));   // memory_op.v(166)
    Mux_4u_16u Mux_597 (.sel({r2_op_inner}), .data({n399, n399, r1[20], 
            a2[20], a1[20], n399, n399, n399, n399, n399, n399, 
            n399, n399, n399, n399, n399}), .o(n598));   // memory_op.v(166)
    Mux_4u_16u Mux_598 (.sel({r2_op_inner}), .data({n400, n400, r1[19], 
            a2[19], a1[19], n400, n400, n400, n400, n400, n400, 
            n400, n400, n400, n400, n400}), .o(n599));   // memory_op.v(166)
    Mux_4u_16u Mux_599 (.sel({r2_op_inner}), .data({n401, n401, r1[18], 
            a2[18], a1[18], n401, n401, n401, n401, n401, n401, 
            n401, n401, n401, n401, n401}), .o(n600));   // memory_op.v(166)
    Mux_4u_16u Mux_600 (.sel({r2_op_inner}), .data({n402, n402, r1[17], 
            a2[17], a1[17], n402, n402, n402, n402, n402, n402, 
            n402, n402, n402, n402, n402}), .o(n601));   // memory_op.v(166)
    Mux_4u_16u Mux_601 (.sel({r2_op_inner}), .data({n403, n403, r1[16], 
            a2[16], a1[16], n403, n403, n403, n403, n403, n403, 
            n403, n403, n403, n403, n403}), .o(n602));   // memory_op.v(166)
    Mux_4u_16u Mux_602 (.sel({r2_op_inner}), .data({n404, n404, r1[15], 
            a2[15], a1[15], n404, n404, n404, n404, n404, n404, 
            n404, n404, n404, n404, n404}), .o(n603));   // memory_op.v(166)
    Mux_4u_16u Mux_603 (.sel({r2_op_inner}), .data({n405, n405, r1[14], 
            a2[14], a1[14], n405, n405, n405, n405, n405, n405, 
            n405, n405, n405, n405, n405}), .o(n604));   // memory_op.v(166)
    Mux_4u_16u Mux_604 (.sel({r2_op_inner}), .data({n406, n406, r1[13], 
            a2[13], a1[13], n406, n406, n406, n406, n406, n406, 
            n406, n406, n406, n406, n406}), .o(n605));   // memory_op.v(166)
    Mux_4u_16u Mux_605 (.sel({r2_op_inner}), .data({n407, n407, r1[12], 
            a2[12], a1[12], n407, n407, n407, n407, n407, n407, 
            n407, n407, n407, n407, n407}), .o(n606));   // memory_op.v(166)
    Mux_4u_16u Mux_606 (.sel({r2_op_inner}), .data({n408, n408, r1[11], 
            a2[11], a1[11], n408, n408, n408, n408, n408, n408, 
            n408, n408, n408, n408, n408}), .o(n607));   // memory_op.v(166)
    Mux_4u_16u Mux_607 (.sel({r2_op_inner}), .data({n409, n409, r1[10], 
            a2[10], a1[10], n409, n409, n409, n409, n409, n409, 
            n409, n409, n409, n409, n409}), .o(n608));   // memory_op.v(166)
    Mux_4u_16u Mux_608 (.sel({r2_op_inner}), .data({n410, n410, r1[9], 
            a2[9], a1[9], n410, n410, n410, n410, n410, n410, 
            n410, n410, n410, n410, n410}), .o(n609));   // memory_op.v(166)
    Mux_4u_16u Mux_609 (.sel({r2_op_inner}), .data({n411, n411, r1[8], 
            a2[8], a1[8], n411, n411, n411, n411, n411, n411, 
            n411, n411, n411, n411, n411}), .o(n610));   // memory_op.v(166)
    Mux_4u_16u Mux_610 (.sel({r2_op_inner}), .data({n412, n412, r1[7], 
            a2[7], a1[7], n412, n412, n412, n412, n412, n412, 
            n412, n412, n412, n412, n412}), .o(n611));   // memory_op.v(166)
    Mux_4u_16u Mux_611 (.sel({r2_op_inner}), .data({n413, n413, r1[6], 
            a2[6], a1[6], n413, n413, n413, n413, n413, n413, 
            n413, n413, n413, n413, n413}), .o(n612));   // memory_op.v(166)
    Mux_4u_16u Mux_612 (.sel({r2_op_inner}), .data({n414, n414, r1[5], 
            a2[5], a1[5], n414, n414, n414, n414, n414, n414, 
            n414, n414, n414, n414, n414}), .o(n613));   // memory_op.v(166)
    Mux_4u_16u Mux_613 (.sel({r2_op_inner}), .data({n415, n415, r1[4], 
            a2[4], a1[4], n415, n415, n415, n415, n415, n415, 
            n415, n415, n415, n415, n415}), .o(n614));   // memory_op.v(166)
    Mux_4u_16u Mux_614 (.sel({r2_op_inner}), .data({n416, n416, r1[3], 
            a2[3], a1[3], n416, n416, n416, n416, n416, n416, 
            n416, n416, n416, n416, n416}), .o(n615));   // memory_op.v(166)
    Mux_4u_16u Mux_615 (.sel({r2_op_inner}), .data({n417, n417, r1[2], 
            a2[2], a1[2], n417, n417, n417, n417, n417, n417, 
            n417, n417, n417, n417, n417}), .o(n616));   // memory_op.v(166)
    Mux_4u_16u Mux_616 (.sel({r2_op_inner}), .data({n418, n418, r1[1], 
            a2[1], a1[1], n418, n418, n418, n418, n418, n418, 
            n418, n418, n418, n418, n418}), .o(n617));   // memory_op.v(166)
    Mux_4u_16u Mux_617 (.sel({r2_op_inner}), .data({n419, n419, r1[0], 
            a2[0], a1[0], n419, n419, n419, n419, n419, n419, 
            n419, n419, n419, n419, n419}), .o(n618));   // memory_op.v(166)
    Mux_4u_16u Mux_618 (.sel({r2_op_inner}), .data({n420, n420, 3'b111, 
            n420, n420, n420, n420, n420, n420, n420, n420, 
            n420, n420, n420}), .o(n619));   // memory_op.v(166)
    Mux_4u_16u Mux_619 (.sel({r2_op_inner}), .data({n421, n421, n421, 
            n421, n421, r1[31], a2[31], a1[31], n421, n421, n421, 
            n421, n421, n421, n421, n421}), .o(n620));   // memory_op.v(166)
    Mux_4u_16u Mux_620 (.sel({r2_op_inner}), .data({n422, n422, n422, 
            n422, n422, r1[30], a2[30], a1[30], n422, n422, n422, 
            n422, n422, n422, n422, n422}), .o(n621));   // memory_op.v(166)
    Mux_4u_16u Mux_621 (.sel({r2_op_inner}), .data({n423, n423, n423, 
            n423, n423, r1[29], a2[29], a1[29], n423, n423, n423, 
            n423, n423, n423, n423, n423}), .o(n622));   // memory_op.v(166)
    Mux_4u_16u Mux_622 (.sel({r2_op_inner}), .data({n424, n424, n424, 
            n424, n424, r1[28], a2[28], a1[28], n424, n424, n424, 
            n424, n424, n424, n424, n424}), .o(n623));   // memory_op.v(166)
    Mux_4u_16u Mux_623 (.sel({r2_op_inner}), .data({n425, n425, n425, 
            n425, n425, r1[27], a2[27], a1[27], n425, n425, n425, 
            n425, n425, n425, n425, n425}), .o(n624));   // memory_op.v(166)
    Mux_4u_16u Mux_624 (.sel({r2_op_inner}), .data({n426, n426, n426, 
            n426, n426, r1[26], a2[26], a1[26], n426, n426, n426, 
            n426, n426, n426, n426, n426}), .o(n625));   // memory_op.v(166)
    Mux_4u_16u Mux_625 (.sel({r2_op_inner}), .data({n427, n427, n427, 
            n427, n427, r1[25], a2[25], a1[25], n427, n427, n427, 
            n427, n427, n427, n427, n427}), .o(n626));   // memory_op.v(166)
    Mux_4u_16u Mux_626 (.sel({r2_op_inner}), .data({n428, n428, n428, 
            n428, n428, r1[24], a2[24], a1[24], n428, n428, n428, 
            n428, n428, n428, n428, n428}), .o(n627));   // memory_op.v(166)
    Mux_4u_16u Mux_627 (.sel({r2_op_inner}), .data({n429, n429, n429, 
            n429, n429, r1[23], a2[23], a1[23], n429, n429, n429, 
            n429, n429, n429, n429, n429}), .o(n628));   // memory_op.v(166)
    Mux_4u_16u Mux_628 (.sel({r2_op_inner}), .data({n430, n430, n430, 
            n430, n430, r1[22], a2[22], a1[22], n430, n430, n430, 
            n430, n430, n430, n430, n430}), .o(n629));   // memory_op.v(166)
    Mux_4u_16u Mux_629 (.sel({r2_op_inner}), .data({n431, n431, n431, 
            n431, n431, r1[21], a2[21], a1[21], n431, n431, n431, 
            n431, n431, n431, n431, n431}), .o(n630));   // memory_op.v(166)
    Mux_4u_16u Mux_630 (.sel({r2_op_inner}), .data({n432, n432, n432, 
            n432, n432, r1[20], a2[20], a1[20], n432, n432, n432, 
            n432, n432, n432, n432, n432}), .o(n631));   // memory_op.v(166)
    Mux_4u_16u Mux_631 (.sel({r2_op_inner}), .data({n433, n433, n433, 
            n433, n433, r1[19], a2[19], a1[19], n433, n433, n433, 
            n433, n433, n433, n433, n433}), .o(n632));   // memory_op.v(166)
    Mux_4u_16u Mux_632 (.sel({r2_op_inner}), .data({n434, n434, n434, 
            n434, n434, r1[18], a2[18], a1[18], n434, n434, n434, 
            n434, n434, n434, n434, n434}), .o(n633));   // memory_op.v(166)
    Mux_4u_16u Mux_633 (.sel({r2_op_inner}), .data({n435, n435, n435, 
            n435, n435, r1[17], a2[17], a1[17], n435, n435, n435, 
            n435, n435, n435, n435, n435}), .o(n634));   // memory_op.v(166)
    Mux_4u_16u Mux_634 (.sel({r2_op_inner}), .data({n436, n436, n436, 
            n436, n436, r1[16], a2[16], a1[16], n436, n436, n436, 
            n436, n436, n436, n436, n436}), .o(n635));   // memory_op.v(166)
    Mux_4u_16u Mux_635 (.sel({r2_op_inner}), .data({n437, n437, n437, 
            n437, n437, r1[15], a2[15], a1[15], n437, n437, n437, 
            n437, n437, n437, n437, n437}), .o(n636));   // memory_op.v(166)
    Mux_4u_16u Mux_636 (.sel({r2_op_inner}), .data({n438, n438, n438, 
            n438, n438, r1[14], a2[14], a1[14], n438, n438, n438, 
            n438, n438, n438, n438, n438}), .o(n637));   // memory_op.v(166)
    Mux_4u_16u Mux_637 (.sel({r2_op_inner}), .data({n439, n439, n439, 
            n439, n439, r1[13], a2[13], a1[13], n439, n439, n439, 
            n439, n439, n439, n439, n439}), .o(n638));   // memory_op.v(166)
    Mux_4u_16u Mux_638 (.sel({r2_op_inner}), .data({n440, n440, n440, 
            n440, n440, r1[12], a2[12], a1[12], n440, n440, n440, 
            n440, n440, n440, n440, n440}), .o(n639));   // memory_op.v(166)
    Mux_4u_16u Mux_639 (.sel({r2_op_inner}), .data({n441, n441, n441, 
            n441, n441, r1[11], a2[11], a1[11], n441, n441, n441, 
            n441, n441, n441, n441, n441}), .o(n640));   // memory_op.v(166)
    Mux_4u_16u Mux_640 (.sel({r2_op_inner}), .data({n442, n442, n442, 
            n442, n442, r1[10], a2[10], a1[10], n442, n442, n442, 
            n442, n442, n442, n442, n442}), .o(n641));   // memory_op.v(166)
    Mux_4u_16u Mux_641 (.sel({r2_op_inner}), .data({n443, n443, n443, 
            n443, n443, r1[9], a2[9], a1[9], n443, n443, n443, 
            n443, n443, n443, n443, n443}), .o(n642));   // memory_op.v(166)
    Mux_4u_16u Mux_642 (.sel({r2_op_inner}), .data({n444, n444, n444, 
            n444, n444, r1[8], a2[8], a1[8], n444, n444, n444, 
            n444, n444, n444, n444, n444}), .o(n643));   // memory_op.v(166)
    Mux_4u_16u Mux_643 (.sel({r2_op_inner}), .data({n445, n445, n445, 
            n445, n445, r1[7], a2[7], a1[7], n445, n445, n445, 
            n445, n445, n445, n445, n445}), .o(n644));   // memory_op.v(166)
    Mux_4u_16u Mux_644 (.sel({r2_op_inner}), .data({n446, n446, n446, 
            n446, n446, r1[6], a2[6], a1[6], n446, n446, n446, 
            n446, n446, n446, n446, n446}), .o(n645));   // memory_op.v(166)
    Mux_4u_16u Mux_645 (.sel({r2_op_inner}), .data({n447, n447, n447, 
            n447, n447, r1[5], a2[5], a1[5], n447, n447, n447, 
            n447, n447, n447, n447, n447}), .o(n646));   // memory_op.v(166)
    Mux_4u_16u Mux_646 (.sel({r2_op_inner}), .data({n448, n448, n448, 
            n448, n448, r1[4], a2[4], a1[4], n448, n448, n448, 
            n448, n448, n448, n448, n448}), .o(n647));   // memory_op.v(166)
    Mux_4u_16u Mux_647 (.sel({r2_op_inner}), .data({n449, n449, n449, 
            n449, n449, r1[3], a2[3], a1[3], n449, n449, n449, 
            n449, n449, n449, n449, n449}), .o(n648));   // memory_op.v(166)
    Mux_4u_16u Mux_648 (.sel({r2_op_inner}), .data({n450, n450, n450, 
            n450, n450, r1[2], a2[2], a1[2], n450, n450, n450, 
            n450, n450, n450, n450, n450}), .o(n649));   // memory_op.v(166)
    Mux_4u_16u Mux_649 (.sel({r2_op_inner}), .data({n451, n451, n451, 
            n451, n451, r1[1], a2[1], a1[1], n451, n451, n451, 
            n451, n451, n451, n451, n451}), .o(n650));   // memory_op.v(166)
    Mux_4u_16u Mux_650 (.sel({r2_op_inner}), .data({n452, n452, n452, 
            n452, n452, r1[0], a2[0], a1[0], n452, n452, n452, 
            n452, n452, n452, n452, n452}), .o(n651));   // memory_op.v(166)
    Mux_4u_16u Mux_651 (.sel({r2_op_inner}), .data({n453, n453, n453, 
            n453, n453, 3'b111, n453, n453, n453, n453, n453, 
            n453, n453, n453}), .o(n652));   // memory_op.v(166)
    Mux_4u_16u Mux_652 (.sel({r2_op_inner}), .data({n454, n454, n454, 
            n454, n454, n454, n454, n454, r2[31], r2[31], r2[31], 
            n454, n454, n454, n454, n454}), .o(n653));   // memory_op.v(166)
    Mux_4u_16u Mux_653 (.sel({r2_op_inner}), .data({n455, n455, n455, 
            n455, n455, n455, n455, n455, r2[30], r2[30], r2[30], 
            n455, n455, n455, n455, n455}), .o(n654));   // memory_op.v(166)
    Mux_4u_16u Mux_654 (.sel({r2_op_inner}), .data({n456, n456, n456, 
            n456, n456, n456, n456, n456, r2[29], r2[29], r2[29], 
            n456, n456, n456, n456, n456}), .o(n655));   // memory_op.v(166)
    Mux_4u_16u Mux_655 (.sel({r2_op_inner}), .data({n457, n457, n457, 
            n457, n457, n457, n457, n457, r2[28], r2[28], r2[28], 
            n457, n457, n457, n457, n457}), .o(n656));   // memory_op.v(166)
    Mux_4u_16u Mux_656 (.sel({r2_op_inner}), .data({n458, n458, n458, 
            n458, n458, n458, n458, n458, r2[27], r2[27], r2[27], 
            n458, n458, n458, n458, n458}), .o(n657));   // memory_op.v(166)
    Mux_4u_16u Mux_657 (.sel({r2_op_inner}), .data({n459, n459, n459, 
            n459, n459, n459, n459, n459, r2[26], r2[26], r2[26], 
            n459, n459, n459, n459, n459}), .o(n658));   // memory_op.v(166)
    Mux_4u_16u Mux_658 (.sel({r2_op_inner}), .data({n460, n460, n460, 
            n460, n460, n460, n460, n460, r2[25], r2[25], r2[25], 
            n460, n460, n460, n460, n460}), .o(n659));   // memory_op.v(166)
    Mux_4u_16u Mux_659 (.sel({r2_op_inner}), .data({n461, n461, n461, 
            n461, n461, n461, n461, n461, r2[24], r2[24], r2[24], 
            n461, n461, n461, n461, n461}), .o(n660));   // memory_op.v(166)
    Mux_4u_16u Mux_660 (.sel({r2_op_inner}), .data({n462, n462, n462, 
            n462, n462, n462, n462, n462, r2[23], r2[23], r2[23], 
            n462, n462, n462, n462, n462}), .o(n661));   // memory_op.v(166)
    Mux_4u_16u Mux_661 (.sel({r2_op_inner}), .data({n463, n463, n463, 
            n463, n463, n463, n463, n463, r2[22], r2[22], r2[22], 
            n463, n463, n463, n463, n463}), .o(n662));   // memory_op.v(166)
    Mux_4u_16u Mux_662 (.sel({r2_op_inner}), .data({n464, n464, n464, 
            n464, n464, n464, n464, n464, r2[21], r2[21], r2[21], 
            n464, n464, n464, n464, n464}), .o(n663));   // memory_op.v(166)
    Mux_4u_16u Mux_663 (.sel({r2_op_inner}), .data({n465, n465, n465, 
            n465, n465, n465, n465, n465, r2[20], r2[20], r2[20], 
            n465, n465, n465, n465, n465}), .o(n664));   // memory_op.v(166)
    Mux_4u_16u Mux_664 (.sel({r2_op_inner}), .data({n466, n466, n466, 
            n466, n466, n466, n466, n466, r2[19], r2[19], r2[19], 
            n466, n466, n466, n466, n466}), .o(n665));   // memory_op.v(166)
    Mux_4u_16u Mux_665 (.sel({r2_op_inner}), .data({n467, n467, n467, 
            n467, n467, n467, n467, n467, r2[18], r2[18], r2[18], 
            n467, n467, n467, n467, n467}), .o(n666));   // memory_op.v(166)
    Mux_4u_16u Mux_666 (.sel({r2_op_inner}), .data({n468, n468, n468, 
            n468, n468, n468, n468, n468, r2[17], r2[17], r2[17], 
            n468, n468, n468, n468, n468}), .o(n667));   // memory_op.v(166)
    Mux_4u_16u Mux_667 (.sel({r2_op_inner}), .data({n469, n469, n469, 
            n469, n469, n469, n469, n469, r2[16], r2[16], r2[16], 
            n469, n469, n469, n469, n469}), .o(n668));   // memory_op.v(166)
    Mux_4u_16u Mux_668 (.sel({r2_op_inner}), .data({n470, n470, n470, 
            n470, n470, n470, n470, n470, r2[15], r2[15], r2[15], 
            n470, n470, n470, n470, n470}), .o(n669));   // memory_op.v(166)
    Mux_4u_16u Mux_669 (.sel({r2_op_inner}), .data({n471, n471, n471, 
            n471, n471, n471, n471, n471, r2[14], r2[14], r2[14], 
            n471, n471, n471, n471, n471}), .o(n670));   // memory_op.v(166)
    Mux_4u_16u Mux_670 (.sel({r2_op_inner}), .data({n472, n472, n472, 
            n472, n472, n472, n472, n472, r2[13], r2[13], r2[13], 
            n472, n472, n472, n472, n472}), .o(n671));   // memory_op.v(166)
    Mux_4u_16u Mux_671 (.sel({r2_op_inner}), .data({n473, n473, n473, 
            n473, n473, n473, n473, n473, r2[12], r2[12], r2[12], 
            n473, n473, n473, n473, n473}), .o(n672));   // memory_op.v(166)
    Mux_4u_16u Mux_672 (.sel({r2_op_inner}), .data({n474, n474, n474, 
            n474, n474, n474, n474, n474, r2[11], r2[11], r2[11], 
            n474, n474, n474, n474, n474}), .o(n673));   // memory_op.v(166)
    Mux_4u_16u Mux_673 (.sel({r2_op_inner}), .data({n475, n475, n475, 
            n475, n475, n475, n475, n475, r2[10], r2[10], r2[10], 
            n475, n475, n475, n475, n475}), .o(n674));   // memory_op.v(166)
    Mux_4u_16u Mux_674 (.sel({r2_op_inner}), .data({n476, n476, n476, 
            n476, n476, n476, n476, n476, r2[9], r2[9], r2[9], 
            n476, n476, n476, n476, n476}), .o(n675));   // memory_op.v(166)
    Mux_4u_16u Mux_675 (.sel({r2_op_inner}), .data({n477, n477, n477, 
            n477, n477, n477, n477, n477, r2[8], r2[8], r2[8], 
            n477, n477, n477, n477, n477}), .o(n676));   // memory_op.v(166)
    Mux_4u_16u Mux_676 (.sel({r2_op_inner}), .data({n478, n478, n478, 
            n478, n478, n478, n478, n478, r2[7], r2[7], r2[7], 
            n478, n478, n478, n478, n478}), .o(n677));   // memory_op.v(166)
    Mux_4u_16u Mux_677 (.sel({r2_op_inner}), .data({n479, n479, n479, 
            n479, n479, n479, n479, n479, r2[6], r2[6], r2[6], 
            n479, n479, n479, n479, n479}), .o(n678));   // memory_op.v(166)
    Mux_4u_16u Mux_678 (.sel({r2_op_inner}), .data({n480, n480, n480, 
            n480, n480, n480, n480, n480, r2[5], r2[5], r2[5], 
            n480, n480, n480, n480, n480}), .o(n679));   // memory_op.v(166)
    Mux_4u_16u Mux_679 (.sel({r2_op_inner}), .data({n481, n481, n481, 
            n481, n481, n481, n481, n481, r2[4], r2[4], r2[4], 
            n481, n481, n481, n481, n481}), .o(n680));   // memory_op.v(166)
    Mux_4u_16u Mux_680 (.sel({r2_op_inner}), .data({n482, n482, n482, 
            n482, n482, n482, n482, n482, r2[3], r2[3], r2[3], 
            n482, n482, n482, n482, n482}), .o(n681));   // memory_op.v(166)
    Mux_4u_16u Mux_681 (.sel({r2_op_inner}), .data({n483, n483, n483, 
            n483, n483, n483, n483, n483, r2[2], r2[2], r2[2], 
            n483, n483, n483, n483, n483}), .o(n682));   // memory_op.v(166)
    Mux_4u_16u Mux_682 (.sel({r2_op_inner}), .data({n484, n484, n484, 
            n484, n484, n484, n484, n484, r2[1], r2[1], r2[1], 
            n484, n484, n484, n484, n484}), .o(n683));   // memory_op.v(166)
    Mux_4u_16u Mux_683 (.sel({r2_op_inner}), .data({n485, n485, n485, 
            n485, n485, n485, n485, n485, r2[0], r2[0], r2[0], 
            n485, n485, n485, n485, n485}), .o(n684));   // memory_op.v(166)
    Mux_4u_16u Mux_684 (.sel({r2_op_inner}), .data({n486, n486, n486, 
            n486, n486, n486, n486, n486, r1[31], a2[31], a1[31], 
            n486, n486, n486, n486, n486}), .o(n685));   // memory_op.v(166)
    Mux_4u_16u Mux_685 (.sel({r2_op_inner}), .data({n487, n487, n487, 
            n487, n487, n487, n487, n487, r1[30], a2[30], a1[30], 
            n487, n487, n487, n487, n487}), .o(n686));   // memory_op.v(166)
    Mux_4u_16u Mux_686 (.sel({r2_op_inner}), .data({n488, n488, n488, 
            n488, n488, n488, n488, n488, r1[29], a2[29], a1[29], 
            n488, n488, n488, n488, n488}), .o(n687));   // memory_op.v(166)
    Mux_4u_16u Mux_687 (.sel({r2_op_inner}), .data({n489, n489, n489, 
            n489, n489, n489, n489, n489, r1[28], a2[28], a1[28], 
            n489, n489, n489, n489, n489}), .o(n688));   // memory_op.v(166)
    Mux_4u_16u Mux_688 (.sel({r2_op_inner}), .data({n490, n490, n490, 
            n490, n490, n490, n490, n490, r1[27], a2[27], a1[27], 
            n490, n490, n490, n490, n490}), .o(n689));   // memory_op.v(166)
    Mux_4u_16u Mux_689 (.sel({r2_op_inner}), .data({n491, n491, n491, 
            n491, n491, n491, n491, n491, r1[26], a2[26], a1[26], 
            n491, n491, n491, n491, n491}), .o(n690));   // memory_op.v(166)
    Mux_4u_16u Mux_690 (.sel({r2_op_inner}), .data({n492, n492, n492, 
            n492, n492, n492, n492, n492, r1[25], a2[25], a1[25], 
            n492, n492, n492, n492, n492}), .o(n691));   // memory_op.v(166)
    Mux_4u_16u Mux_691 (.sel({r2_op_inner}), .data({n493, n493, n493, 
            n493, n493, n493, n493, n493, r1[24], a2[24], a1[24], 
            n493, n493, n493, n493, n493}), .o(n692));   // memory_op.v(166)
    Mux_4u_16u Mux_692 (.sel({r2_op_inner}), .data({n494, n494, n494, 
            n494, n494, n494, n494, n494, r1[23], a2[23], a1[23], 
            n494, n494, n494, n494, n494}), .o(n693));   // memory_op.v(166)
    Mux_4u_16u Mux_693 (.sel({r2_op_inner}), .data({n495, n495, n495, 
            n495, n495, n495, n495, n495, r1[22], a2[22], a1[22], 
            n495, n495, n495, n495, n495}), .o(n694));   // memory_op.v(166)
    Mux_4u_16u Mux_694 (.sel({r2_op_inner}), .data({n496, n496, n496, 
            n496, n496, n496, n496, n496, r1[21], a2[21], a1[21], 
            n496, n496, n496, n496, n496}), .o(n695));   // memory_op.v(166)
    Mux_4u_16u Mux_695 (.sel({r2_op_inner}), .data({n497, n497, n497, 
            n497, n497, n497, n497, n497, r1[20], a2[20], a1[20], 
            n497, n497, n497, n497, n497}), .o(n696));   // memory_op.v(166)
    Mux_4u_16u Mux_696 (.sel({r2_op_inner}), .data({n498, n498, n498, 
            n498, n498, n498, n498, n498, r1[19], a2[19], a1[19], 
            n498, n498, n498, n498, n498}), .o(n697));   // memory_op.v(166)
    Mux_4u_16u Mux_697 (.sel({r2_op_inner}), .data({n499, n499, n499, 
            n499, n499, n499, n499, n499, r1[18], a2[18], a1[18], 
            n499, n499, n499, n499, n499}), .o(n698));   // memory_op.v(166)
    Mux_4u_16u Mux_698 (.sel({r2_op_inner}), .data({n500, n500, n500, 
            n500, n500, n500, n500, n500, r1[17], a2[17], a1[17], 
            n500, n500, n500, n500, n500}), .o(n699));   // memory_op.v(166)
    Mux_4u_16u Mux_699 (.sel({r2_op_inner}), .data({n501, n501, n501, 
            n501, n501, n501, n501, n501, r1[16], a2[16], a1[16], 
            n501, n501, n501, n501, n501}), .o(n700));   // memory_op.v(166)
    Mux_4u_16u Mux_700 (.sel({r2_op_inner}), .data({n502, n502, n502, 
            n502, n502, n502, n502, n502, r1[15], a2[15], a1[15], 
            n502, n502, n502, n502, n502}), .o(n701));   // memory_op.v(166)
    Mux_4u_16u Mux_701 (.sel({r2_op_inner}), .data({n503, n503, n503, 
            n503, n503, n503, n503, n503, r1[14], a2[14], a1[14], 
            n503, n503, n503, n503, n503}), .o(n702));   // memory_op.v(166)
    Mux_4u_16u Mux_702 (.sel({r2_op_inner}), .data({n504, n504, n504, 
            n504, n504, n504, n504, n504, r1[13], a2[13], a1[13], 
            n504, n504, n504, n504, n504}), .o(n703));   // memory_op.v(166)
    Mux_4u_16u Mux_703 (.sel({r2_op_inner}), .data({n505, n505, n505, 
            n505, n505, n505, n505, n505, r1[12], a2[12], a1[12], 
            n505, n505, n505, n505, n505}), .o(n704));   // memory_op.v(166)
    Mux_4u_16u Mux_704 (.sel({r2_op_inner}), .data({n506, n506, n506, 
            n506, n506, n506, n506, n506, r1[11], a2[11], a1[11], 
            n506, n506, n506, n506, n506}), .o(n705));   // memory_op.v(166)
    Mux_4u_16u Mux_705 (.sel({r2_op_inner}), .data({n507, n507, n507, 
            n507, n507, n507, n507, n507, r1[10], a2[10], a1[10], 
            n507, n507, n507, n507, n507}), .o(n706));   // memory_op.v(166)
    Mux_4u_16u Mux_706 (.sel({r2_op_inner}), .data({n508, n508, n508, 
            n508, n508, n508, n508, n508, r1[9], a2[9], a1[9], 
            n508, n508, n508, n508, n508}), .o(n707));   // memory_op.v(166)
    Mux_4u_16u Mux_707 (.sel({r2_op_inner}), .data({n509, n509, n509, 
            n509, n509, n509, n509, n509, r1[8], a2[8], a1[8], 
            n509, n509, n509, n509, n509}), .o(n708));   // memory_op.v(166)
    Mux_4u_16u Mux_708 (.sel({r2_op_inner}), .data({n510, n510, n510, 
            n510, n510, n510, n510, n510, r1[7], a2[7], a1[7], 
            n510, n510, n510, n510, n510}), .o(n709));   // memory_op.v(166)
    Mux_4u_16u Mux_709 (.sel({r2_op_inner}), .data({n511, n511, n511, 
            n511, n511, n511, n511, n511, r1[6], a2[6], a1[6], 
            n511, n511, n511, n511, n511}), .o(n710));   // memory_op.v(166)
    Mux_4u_16u Mux_710 (.sel({r2_op_inner}), .data({n512, n512, n512, 
            n512, n512, n512, n512, n512, r1[5], a2[5], a1[5], 
            n512, n512, n512, n512, n512}), .o(n711));   // memory_op.v(166)
    Mux_4u_16u Mux_711 (.sel({r2_op_inner}), .data({n513, n513, n513, 
            n513, n513, n513, n513, n513, r1[4], a2[4], a1[4], 
            n513, n513, n513, n513, n513}), .o(n712));   // memory_op.v(166)
    Mux_4u_16u Mux_712 (.sel({r2_op_inner}), .data({n514, n514, n514, 
            n514, n514, n514, n514, n514, r1[3], a2[3], a1[3], 
            n514, n514, n514, n514, n514}), .o(n713));   // memory_op.v(166)
    Mux_4u_16u Mux_713 (.sel({r2_op_inner}), .data({n515, n515, n515, 
            n515, n515, n515, n515, n515, r1[2], a2[2], a1[2], 
            n515, n515, n515, n515, n515}), .o(n714));   // memory_op.v(166)
    Mux_4u_16u Mux_714 (.sel({r2_op_inner}), .data({n516, n516, n516, 
            n516, n516, n516, n516, n516, r1[1], a2[1], a1[1], 
            n516, n516, n516, n516, n516}), .o(n715));   // memory_op.v(166)
    Mux_4u_16u Mux_715 (.sel({r2_op_inner}), .data({n517, n517, n517, 
            n517, n517, n517, n517, n517, r1[0], a2[0], a1[0], 
            n517, n517, n517, n517, n517}), .o(n716));   // memory_op.v(166)
    Mux_4u_16u Mux_716 (.sel({r2_op_inner}), .data({n518, n518, n518, 
            n518, n518, n518, n518, n518, 3'b111, n518, n518, 
            n518, n518, n518}), .o(n717));   // memory_op.v(166)
    Mux_4u_16u Mux_717 (.sel({r2_op_inner}), .data({n519, n519, n519, 
            n519, n519, n519, n519, n519, n519, n519, n519, 
            r1[31], a2[31], a1[31], n519, n519}), .o(n718));   // memory_op.v(166)
    Mux_4u_16u Mux_718 (.sel({r2_op_inner}), .data({n520, n520, n520, 
            n520, n520, n520, n520, n520, n520, n520, n520, 
            r1[30], a2[30], a1[30], n520, n520}), .o(n719));   // memory_op.v(166)
    Mux_4u_16u Mux_719 (.sel({r2_op_inner}), .data({n521, n521, n521, 
            n521, n521, n521, n521, n521, n521, n521, n521, 
            r1[29], a2[29], a1[29], n521, n521}), .o(n720));   // memory_op.v(166)
    Mux_4u_16u Mux_720 (.sel({r2_op_inner}), .data({n522, n522, n522, 
            n522, n522, n522, n522, n522, n522, n522, n522, 
            r1[28], a2[28], a1[28], n522, n522}), .o(n721));   // memory_op.v(166)
    Mux_4u_16u Mux_721 (.sel({r2_op_inner}), .data({n523, n523, n523, 
            n523, n523, n523, n523, n523, n523, n523, n523, 
            r1[27], a2[27], a1[27], n523, n523}), .o(n722));   // memory_op.v(166)
    Mux_4u_16u Mux_722 (.sel({r2_op_inner}), .data({n524, n524, n524, 
            n524, n524, n524, n524, n524, n524, n524, n524, 
            r1[26], a2[26], a1[26], n524, n524}), .o(n723));   // memory_op.v(166)
    Mux_4u_16u Mux_723 (.sel({r2_op_inner}), .data({n525, n525, n525, 
            n525, n525, n525, n525, n525, n525, n525, n525, 
            r1[25], a2[25], a1[25], n525, n525}), .o(n724));   // memory_op.v(166)
    Mux_4u_16u Mux_724 (.sel({r2_op_inner}), .data({n526, n526, n526, 
            n526, n526, n526, n526, n526, n526, n526, n526, 
            r1[24], a2[24], a1[24], n526, n526}), .o(n725));   // memory_op.v(166)
    Mux_4u_16u Mux_725 (.sel({r2_op_inner}), .data({n527, n527, n527, 
            n527, n527, n527, n527, n527, n527, n527, n527, 
            r1[23], a2[23], a1[23], n527, n527}), .o(n726));   // memory_op.v(166)
    Mux_4u_16u Mux_726 (.sel({r2_op_inner}), .data({n528, n528, n528, 
            n528, n528, n528, n528, n528, n528, n528, n528, 
            r1[22], a2[22], a1[22], n528, n528}), .o(n727));   // memory_op.v(166)
    Mux_4u_16u Mux_727 (.sel({r2_op_inner}), .data({n529, n529, n529, 
            n529, n529, n529, n529, n529, n529, n529, n529, 
            r1[21], a2[21], a1[21], n529, n529}), .o(n728));   // memory_op.v(166)
    Mux_4u_16u Mux_728 (.sel({r2_op_inner}), .data({n530, n530, n530, 
            n530, n530, n530, n530, n530, n530, n530, n530, 
            r1[20], a2[20], a1[20], n530, n530}), .o(n729));   // memory_op.v(166)
    Mux_4u_16u Mux_729 (.sel({r2_op_inner}), .data({n531, n531, n531, 
            n531, n531, n531, n531, n531, n531, n531, n531, 
            r1[19], a2[19], a1[19], n531, n531}), .o(n730));   // memory_op.v(166)
    Mux_4u_16u Mux_730 (.sel({r2_op_inner}), .data({n532, n532, n532, 
            n532, n532, n532, n532, n532, n532, n532, n532, 
            r1[18], a2[18], a1[18], n532, n532}), .o(n731));   // memory_op.v(166)
    Mux_4u_16u Mux_731 (.sel({r2_op_inner}), .data({n533, n533, n533, 
            n533, n533, n533, n533, n533, n533, n533, n533, 
            r1[17], a2[17], a1[17], n533, n533}), .o(n732));   // memory_op.v(166)
    Mux_4u_16u Mux_732 (.sel({r2_op_inner}), .data({n534, n534, n534, 
            n534, n534, n534, n534, n534, n534, n534, n534, 
            r1[16], a2[16], a1[16], n534, n534}), .o(n733));   // memory_op.v(166)
    Mux_4u_16u Mux_733 (.sel({r2_op_inner}), .data({n535, n535, n535, 
            n535, n535, n535, n535, n535, n535, n535, n535, 
            r1[15], a2[15], a1[15], n535, n535}), .o(n734));   // memory_op.v(166)
    Mux_4u_16u Mux_734 (.sel({r2_op_inner}), .data({n536, n536, n536, 
            n536, n536, n536, n536, n536, n536, n536, n536, 
            r1[14], a2[14], a1[14], n536, n536}), .o(n735));   // memory_op.v(166)
    Mux_4u_16u Mux_735 (.sel({r2_op_inner}), .data({n537, n537, n537, 
            n537, n537, n537, n537, n537, n537, n537, n537, 
            r1[13], a2[13], a1[13], n537, n537}), .o(n736));   // memory_op.v(166)
    Mux_4u_16u Mux_736 (.sel({r2_op_inner}), .data({n538, n538, n538, 
            n538, n538, n538, n538, n538, n538, n538, n538, 
            r1[12], a2[12], a1[12], n538, n538}), .o(n737));   // memory_op.v(166)
    Mux_4u_16u Mux_737 (.sel({r2_op_inner}), .data({n539, n539, n539, 
            n539, n539, n539, n539, n539, n539, n539, n539, 
            r1[11], a2[11], a1[11], n539, n539}), .o(n738));   // memory_op.v(166)
    Mux_4u_16u Mux_738 (.sel({r2_op_inner}), .data({n540, n540, n540, 
            n540, n540, n540, n540, n540, n540, n540, n540, 
            r1[10], a2[10], a1[10], n540, n540}), .o(n739));   // memory_op.v(166)
    Mux_4u_16u Mux_739 (.sel({r2_op_inner}), .data({n541, n541, n541, 
            n541, n541, n541, n541, n541, n541, n541, n541, 
            r1[9], a2[9], a1[9], n541, n541}), .o(n740));   // memory_op.v(166)
    Mux_4u_16u Mux_740 (.sel({r2_op_inner}), .data({n542, n542, n542, 
            n542, n542, n542, n542, n542, n542, n542, n542, 
            r1[8], a2[8], a1[8], n542, n542}), .o(n741));   // memory_op.v(166)
    Mux_4u_16u Mux_741 (.sel({r2_op_inner}), .data({n543, n543, n543, 
            n543, n543, n543, n543, n543, n543, n543, n543, 
            r1[7], a2[7], a1[7], n543, n543}), .o(n742));   // memory_op.v(166)
    Mux_4u_16u Mux_742 (.sel({r2_op_inner}), .data({n544, n544, n544, 
            n544, n544, n544, n544, n544, n544, n544, n544, 
            r1[6], a2[6], a1[6], n544, n544}), .o(n743));   // memory_op.v(166)
    Mux_4u_16u Mux_743 (.sel({r2_op_inner}), .data({n545, n545, n545, 
            n545, n545, n545, n545, n545, n545, n545, n545, 
            r1[5], a2[5], a1[5], n545, n545}), .o(n744));   // memory_op.v(166)
    Mux_4u_16u Mux_744 (.sel({r2_op_inner}), .data({n546, n546, n546, 
            n546, n546, n546, n546, n546, n546, n546, n546, 
            r1[4], a2[4], a1[4], n546, n546}), .o(n745));   // memory_op.v(166)
    Mux_4u_16u Mux_745 (.sel({r2_op_inner}), .data({n547, n547, n547, 
            n547, n547, n547, n547, n547, n547, n547, n547, 
            r1[3], a2[3], a1[3], n547, n547}), .o(n746));   // memory_op.v(166)
    Mux_4u_16u Mux_746 (.sel({r2_op_inner}), .data({n548, n548, n548, 
            n548, n548, n548, n548, n548, n548, n548, n548, 
            r1[2], a2[2], a1[2], n548, n548}), .o(n747));   // memory_op.v(166)
    Mux_4u_16u Mux_747 (.sel({r2_op_inner}), .data({n549, n549, n549, 
            n549, n549, n549, n549, n549, n549, n549, n549, 
            r1[1], a2[1], a1[1], n549, n549}), .o(n748));   // memory_op.v(166)
    Mux_4u_16u Mux_748 (.sel({r2_op_inner}), .data({n550, n550, n550, 
            n550, n550, n550, n550, n550, n550, n550, n550, 
            r1[0], a2[0], a1[0], n550, n550}), .o(n749));   // memory_op.v(166)
    Mux_4u_16u Mux_749 (.sel({r2_op_inner}), .data({n551, n551, n551, 
            n551, n551, n551, n551, n551, n551, n551, n551, 
            3'b111, n551, n551}), .o(n750));   // memory_op.v(166)
    VERIFIC_DFFRS i752 (.d(n686), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[30]));   // memory_op.v(69)
    VERIFIC_DFFRS i753 (.d(n687), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[29]));   // memory_op.v(69)
    VERIFIC_DFFRS i754 (.d(n688), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[28]));   // memory_op.v(69)
    VERIFIC_DFFRS i755 (.d(n689), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[27]));   // memory_op.v(69)
    VERIFIC_DFFRS i756 (.d(n690), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[26]));   // memory_op.v(69)
    VERIFIC_DFFRS i757 (.d(n691), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[25]));   // memory_op.v(69)
    VERIFIC_DFFRS i758 (.d(n692), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[24]));   // memory_op.v(69)
    VERIFIC_DFFRS i759 (.d(n693), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[23]));   // memory_op.v(69)
    VERIFIC_DFFRS i760 (.d(n694), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[22]));   // memory_op.v(69)
    VERIFIC_DFFRS i761 (.d(n695), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[21]));   // memory_op.v(69)
    VERIFIC_DFFRS i762 (.d(n696), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[20]));   // memory_op.v(69)
    VERIFIC_DFFRS i763 (.d(n697), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[19]));   // memory_op.v(69)
    VERIFIC_DFFRS i764 (.d(n698), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[18]));   // memory_op.v(69)
    VERIFIC_DFFRS i765 (.d(n699), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[17]));   // memory_op.v(69)
    VERIFIC_DFFRS i766 (.d(n700), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[16]));   // memory_op.v(69)
    VERIFIC_DFFRS i767 (.d(n701), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[15]));   // memory_op.v(69)
    VERIFIC_DFFRS i768 (.d(n702), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[14]));   // memory_op.v(69)
    VERIFIC_DFFRS i769 (.d(n703), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[13]));   // memory_op.v(69)
    VERIFIC_DFFRS i770 (.d(n704), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[12]));   // memory_op.v(69)
    VERIFIC_DFFRS i771 (.d(n705), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[11]));   // memory_op.v(69)
    VERIFIC_DFFRS i772 (.d(n706), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[10]));   // memory_op.v(69)
    VERIFIC_DFFRS i773 (.d(n707), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[9]));   // memory_op.v(69)
    VERIFIC_DFFRS i774 (.d(n708), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[8]));   // memory_op.v(69)
    VERIFIC_DFFRS i775 (.d(n709), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[7]));   // memory_op.v(69)
    VERIFIC_DFFRS i776 (.d(n710), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[6]));   // memory_op.v(69)
    VERIFIC_DFFRS i777 (.d(n711), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[5]));   // memory_op.v(69)
    VERIFIC_DFFRS i778 (.d(n712), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[4]));   // memory_op.v(69)
    VERIFIC_DFFRS i779 (.d(n713), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[3]));   // memory_op.v(69)
    VERIFIC_DFFRS i780 (.d(n714), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[2]));   // memory_op.v(69)
    VERIFIC_DFFRS i781 (.d(n715), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[1]));   // memory_op.v(69)
    VERIFIC_DFFRS i782 (.d(n716), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[0]));   // memory_op.v(69)
    VERIFIC_DFFRS i783 (.d(n718), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[31]));   // memory_op.v(69)
    VERIFIC_DFFRS i784 (.d(n719), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[30]));   // memory_op.v(69)
    VERIFIC_DFFRS i785 (.d(n720), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[29]));   // memory_op.v(69)
    VERIFIC_DFFRS i786 (.d(n721), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[28]));   // memory_op.v(69)
    VERIFIC_DFFRS i787 (.d(n722), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[27]));   // memory_op.v(69)
    VERIFIC_DFFRS i788 (.d(n723), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[26]));   // memory_op.v(69)
    VERIFIC_DFFRS i789 (.d(n724), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[25]));   // memory_op.v(69)
    VERIFIC_DFFRS i790 (.d(n725), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[24]));   // memory_op.v(69)
    VERIFIC_DFFRS i791 (.d(n726), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[23]));   // memory_op.v(69)
    VERIFIC_DFFRS i792 (.d(n727), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[22]));   // memory_op.v(69)
    VERIFIC_DFFRS i793 (.d(n728), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[21]));   // memory_op.v(69)
    VERIFIC_DFFRS i794 (.d(n729), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[20]));   // memory_op.v(69)
    VERIFIC_DFFRS i795 (.d(n730), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[19]));   // memory_op.v(69)
    VERIFIC_DFFRS i796 (.d(n731), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[18]));   // memory_op.v(69)
    VERIFIC_DFFRS i797 (.d(n732), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[17]));   // memory_op.v(69)
    VERIFIC_DFFRS i798 (.d(n733), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[16]));   // memory_op.v(69)
    VERIFIC_DFFRS i799 (.d(n734), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[15]));   // memory_op.v(69)
    VERIFIC_DFFRS i800 (.d(n735), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[14]));   // memory_op.v(69)
    VERIFIC_DFFRS i801 (.d(n736), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[13]));   // memory_op.v(69)
    VERIFIC_DFFRS i802 (.d(n737), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[12]));   // memory_op.v(69)
    VERIFIC_DFFRS i803 (.d(n738), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[11]));   // memory_op.v(69)
    VERIFIC_DFFRS i804 (.d(n739), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[10]));   // memory_op.v(69)
    VERIFIC_DFFRS i805 (.d(n740), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[9]));   // memory_op.v(69)
    VERIFIC_DFFRS i806 (.d(n741), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[8]));   // memory_op.v(69)
    VERIFIC_DFFRS i807 (.d(n742), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[7]));   // memory_op.v(69)
    VERIFIC_DFFRS i808 (.d(n743), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[6]));   // memory_op.v(69)
    VERIFIC_DFFRS i809 (.d(n744), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[5]));   // memory_op.v(69)
    VERIFIC_DFFRS i810 (.d(n745), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[4]));   // memory_op.v(69)
    VERIFIC_DFFRS i811 (.d(n746), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[3]));   // memory_op.v(69)
    VERIFIC_DFFRS i812 (.d(n747), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[2]));   // memory_op.v(69)
    VERIFIC_DFFRS i813 (.d(n748), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[1]));   // memory_op.v(69)
    VERIFIC_DFFRS i814 (.d(n749), .clk(clk), .s(1'b0), .r(rst), .q(ram_r_addr[0]));   // memory_op.v(69)
    VERIFIC_DFFRS i815 (.d(n587), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[31]));   // memory_op.v(69)
    VERIFIC_DFFRS i816 (.d(n588), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[30]));   // memory_op.v(69)
    VERIFIC_DFFRS i817 (.d(n589), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[29]));   // memory_op.v(69)
    VERIFIC_DFFRS i818 (.d(n590), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[28]));   // memory_op.v(69)
    VERIFIC_DFFRS i819 (.d(n591), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[27]));   // memory_op.v(69)
    VERIFIC_DFFRS i820 (.d(n592), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[26]));   // memory_op.v(69)
    VERIFIC_DFFRS i821 (.d(n593), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[25]));   // memory_op.v(69)
    VERIFIC_DFFRS i822 (.d(n594), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[24]));   // memory_op.v(69)
    VERIFIC_DFFRS i823 (.d(n595), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[23]));   // memory_op.v(69)
    VERIFIC_DFFRS i824 (.d(n596), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[22]));   // memory_op.v(69)
    VERIFIC_DFFRS i825 (.d(n597), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[21]));   // memory_op.v(69)
    VERIFIC_DFFRS i826 (.d(n598), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[20]));   // memory_op.v(69)
    VERIFIC_DFFRS i827 (.d(n599), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[19]));   // memory_op.v(69)
    VERIFIC_DFFRS i828 (.d(n600), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[18]));   // memory_op.v(69)
    VERIFIC_DFFRS i829 (.d(n601), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[17]));   // memory_op.v(69)
    VERIFIC_DFFRS i830 (.d(n602), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[16]));   // memory_op.v(69)
    VERIFIC_DFFRS i831 (.d(n603), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[15]));   // memory_op.v(69)
    VERIFIC_DFFRS i832 (.d(n604), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[14]));   // memory_op.v(69)
    VERIFIC_DFFRS i833 (.d(n605), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[13]));   // memory_op.v(69)
    VERIFIC_DFFRS i834 (.d(n606), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[12]));   // memory_op.v(69)
    VERIFIC_DFFRS i835 (.d(n607), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[11]));   // memory_op.v(69)
    VERIFIC_DFFRS i836 (.d(n608), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[10]));   // memory_op.v(69)
    VERIFIC_DFFRS i837 (.d(n609), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[9]));   // memory_op.v(69)
    VERIFIC_DFFRS i838 (.d(n610), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[8]));   // memory_op.v(69)
    VERIFIC_DFFRS i839 (.d(n611), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[7]));   // memory_op.v(69)
    VERIFIC_DFFRS i840 (.d(n612), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[6]));   // memory_op.v(69)
    VERIFIC_DFFRS i841 (.d(n613), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[5]));   // memory_op.v(69)
    VERIFIC_DFFRS i842 (.d(n614), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[4]));   // memory_op.v(69)
    VERIFIC_DFFRS i843 (.d(n615), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[3]));   // memory_op.v(69)
    VERIFIC_DFFRS i844 (.d(n616), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[2]));   // memory_op.v(69)
    VERIFIC_DFFRS i845 (.d(n617), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[1]));   // memory_op.v(69)
    VERIFIC_DFFRS i846 (.d(n618), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_addr[0]));   // memory_op.v(69)
    VERIFIC_DFFRS i847 (.d(n620), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[31]));   // memory_op.v(69)
    VERIFIC_DFFRS i848 (.d(n621), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[30]));   // memory_op.v(69)
    VERIFIC_DFFRS i849 (.d(n622), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[29]));   // memory_op.v(69)
    VERIFIC_DFFRS i850 (.d(n623), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[28]));   // memory_op.v(69)
    VERIFIC_DFFRS i851 (.d(n624), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[27]));   // memory_op.v(69)
    VERIFIC_DFFRS i852 (.d(n625), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[26]));   // memory_op.v(69)
    VERIFIC_DFFRS i853 (.d(n626), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[25]));   // memory_op.v(69)
    VERIFIC_DFFRS i854 (.d(n627), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[24]));   // memory_op.v(69)
    VERIFIC_DFFRS i855 (.d(n628), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[23]));   // memory_op.v(69)
    VERIFIC_DFFRS i856 (.d(n629), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[22]));   // memory_op.v(69)
    VERIFIC_DFFRS i857 (.d(n630), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[21]));   // memory_op.v(69)
    VERIFIC_DFFRS i858 (.d(n631), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[20]));   // memory_op.v(69)
    VERIFIC_DFFRS i859 (.d(n632), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[19]));   // memory_op.v(69)
    VERIFIC_DFFRS i860 (.d(n633), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[18]));   // memory_op.v(69)
    VERIFIC_DFFRS i861 (.d(n634), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[17]));   // memory_op.v(69)
    VERIFIC_DFFRS i862 (.d(n635), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[16]));   // memory_op.v(69)
    VERIFIC_DFFRS i863 (.d(n636), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[15]));   // memory_op.v(69)
    VERIFIC_DFFRS i864 (.d(n637), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[14]));   // memory_op.v(69)
    VERIFIC_DFFRS i865 (.d(n638), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[13]));   // memory_op.v(69)
    VERIFIC_DFFRS i866 (.d(n639), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[12]));   // memory_op.v(69)
    VERIFIC_DFFRS i867 (.d(n640), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[11]));   // memory_op.v(69)
    VERIFIC_DFFRS i868 (.d(n641), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[10]));   // memory_op.v(69)
    VERIFIC_DFFRS i869 (.d(n642), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[9]));   // memory_op.v(69)
    VERIFIC_DFFRS i870 (.d(n643), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[8]));   // memory_op.v(69)
    VERIFIC_DFFRS i871 (.d(n644), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[7]));   // memory_op.v(69)
    VERIFIC_DFFRS i872 (.d(n645), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[6]));   // memory_op.v(69)
    VERIFIC_DFFRS i873 (.d(n646), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[5]));   // memory_op.v(69)
    VERIFIC_DFFRS i874 (.d(n647), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[4]));   // memory_op.v(69)
    VERIFIC_DFFRS i875 (.d(n648), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[3]));   // memory_op.v(69)
    VERIFIC_DFFRS i876 (.d(n649), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[2]));   // memory_op.v(69)
    VERIFIC_DFFRS i877 (.d(n650), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[1]));   // memory_op.v(69)
    VERIFIC_DFFRS i878 (.d(n651), .clk(clk), .s(1'b0), .r(rst), .q(sys_r_addr[0]));   // memory_op.v(69)
    VERIFIC_DFFRS i879 (.d(n653), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[31]));   // memory_op.v(69)
    VERIFIC_DFFRS i880 (.d(n654), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[30]));   // memory_op.v(69)
    VERIFIC_DFFRS i881 (.d(n655), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[29]));   // memory_op.v(69)
    VERIFIC_DFFRS i882 (.d(n656), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[28]));   // memory_op.v(69)
    VERIFIC_DFFRS i883 (.d(n657), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[27]));   // memory_op.v(69)
    VERIFIC_DFFRS i884 (.d(n658), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[26]));   // memory_op.v(69)
    VERIFIC_DFFRS i885 (.d(n659), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[25]));   // memory_op.v(69)
    VERIFIC_DFFRS i886 (.d(n660), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[24]));   // memory_op.v(69)
    VERIFIC_DFFRS i887 (.d(n661), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[23]));   // memory_op.v(69)
    VERIFIC_DFFRS i888 (.d(n662), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[22]));   // memory_op.v(69)
    VERIFIC_DFFRS i889 (.d(n663), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[21]));   // memory_op.v(69)
    VERIFIC_DFFRS i890 (.d(n664), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[20]));   // memory_op.v(69)
    VERIFIC_DFFRS i891 (.d(n665), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[19]));   // memory_op.v(69)
    VERIFIC_DFFRS i892 (.d(n666), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[18]));   // memory_op.v(69)
    VERIFIC_DFFRS i893 (.d(n667), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[17]));   // memory_op.v(69)
    VERIFIC_DFFRS i894 (.d(n668), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[16]));   // memory_op.v(69)
    VERIFIC_DFFRS i895 (.d(n669), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[15]));   // memory_op.v(69)
    VERIFIC_DFFRS i896 (.d(n670), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[14]));   // memory_op.v(69)
    VERIFIC_DFFRS i897 (.d(n671), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[13]));   // memory_op.v(69)
    VERIFIC_DFFRS i898 (.d(n672), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[12]));   // memory_op.v(69)
    VERIFIC_DFFRS i899 (.d(n673), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[11]));   // memory_op.v(69)
    VERIFIC_DFFRS i900 (.d(n674), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[10]));   // memory_op.v(69)
    VERIFIC_DFFRS i901 (.d(n675), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[9]));   // memory_op.v(69)
    VERIFIC_DFFRS i902 (.d(n676), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[8]));   // memory_op.v(69)
    VERIFIC_DFFRS i903 (.d(n677), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[7]));   // memory_op.v(69)
    VERIFIC_DFFRS i904 (.d(n678), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[6]));   // memory_op.v(69)
    VERIFIC_DFFRS i905 (.d(n679), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[5]));   // memory_op.v(69)
    VERIFIC_DFFRS i906 (.d(n680), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[4]));   // memory_op.v(69)
    VERIFIC_DFFRS i907 (.d(n681), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[3]));   // memory_op.v(69)
    VERIFIC_DFFRS i908 (.d(n682), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[2]));   // memory_op.v(69)
    VERIFIC_DFFRS i909 (.d(n683), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[1]));   // memory_op.v(69)
    VERIFIC_DFFRS i910 (.d(n684), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_line[0]));   // memory_op.v(69)
    VERIFIC_DFFRS i911 (.d(n555), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[31]));   // memory_op.v(69)
    VERIFIC_DFFRS i912 (.d(n556), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[30]));   // memory_op.v(69)
    VERIFIC_DFFRS i913 (.d(n557), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[29]));   // memory_op.v(69)
    VERIFIC_DFFRS i914 (.d(n558), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[28]));   // memory_op.v(69)
    VERIFIC_DFFRS i915 (.d(n559), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[27]));   // memory_op.v(69)
    VERIFIC_DFFRS i916 (.d(n560), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[26]));   // memory_op.v(69)
    VERIFIC_DFFRS i917 (.d(n561), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[25]));   // memory_op.v(69)
    VERIFIC_DFFRS i918 (.d(n562), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[24]));   // memory_op.v(69)
    VERIFIC_DFFRS i919 (.d(n563), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[23]));   // memory_op.v(69)
    VERIFIC_DFFRS i920 (.d(n564), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[22]));   // memory_op.v(69)
    VERIFIC_DFFRS i921 (.d(n565), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[21]));   // memory_op.v(69)
    VERIFIC_DFFRS i922 (.d(n566), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[20]));   // memory_op.v(69)
    VERIFIC_DFFRS i923 (.d(n567), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[19]));   // memory_op.v(69)
    VERIFIC_DFFRS i924 (.d(n568), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[18]));   // memory_op.v(69)
    VERIFIC_DFFRS i925 (.d(n569), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[17]));   // memory_op.v(69)
    VERIFIC_DFFRS i926 (.d(n570), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[16]));   // memory_op.v(69)
    VERIFIC_DFFRS i927 (.d(n571), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[15]));   // memory_op.v(69)
    VERIFIC_DFFRS i928 (.d(n572), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[14]));   // memory_op.v(69)
    VERIFIC_DFFRS i929 (.d(n573), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[13]));   // memory_op.v(69)
    VERIFIC_DFFRS i930 (.d(n574), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[12]));   // memory_op.v(69)
    VERIFIC_DFFRS i931 (.d(n575), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[11]));   // memory_op.v(69)
    VERIFIC_DFFRS i932 (.d(n576), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[10]));   // memory_op.v(69)
    VERIFIC_DFFRS i933 (.d(n577), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[9]));   // memory_op.v(69)
    VERIFIC_DFFRS i934 (.d(n578), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[8]));   // memory_op.v(69)
    VERIFIC_DFFRS i935 (.d(n579), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[7]));   // memory_op.v(69)
    VERIFIC_DFFRS i936 (.d(n580), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[6]));   // memory_op.v(69)
    VERIFIC_DFFRS i937 (.d(n581), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[5]));   // memory_op.v(69)
    VERIFIC_DFFRS i938 (.d(n582), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[4]));   // memory_op.v(69)
    VERIFIC_DFFRS i939 (.d(n583), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[3]));   // memory_op.v(69)
    VERIFIC_DFFRS i940 (.d(n584), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[2]));   // memory_op.v(69)
    VERIFIC_DFFRS i941 (.d(n585), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[1]));   // memory_op.v(69)
    VERIFIC_DFFRS i942 (.d(n586), .clk(clk), .s(1'b0), .r(rst), .q(sys_w_line[0]));   // memory_op.v(69)
    VERIFIC_DFFRS i943 (.d(n717), .clk(clk), .s(1'b0), .r(rst), .q(ram_w));   // memory_op.v(69)
    VERIFIC_DFFRS i944 (.d(n750), .clk(clk), .s(1'b0), .r(rst), .q(ram_r));   // memory_op.v(69)
    VERIFIC_DFFRS i945 (.d(n652), .clk(clk), .s(1'b0), .r(rst), .q(sys_r));   // memory_op.v(69)
    VERIFIC_DFFRS i946 (.d(n619), .clk(clk), .s(1'b0), .r(rst), .q(sys_w));   // memory_op.v(69)
    VERIFIC_DFFRS i947 (.d(n353), .clk(clk), .s(1'b0), .r(rst), .q(m1_select[2]));   // memory_op.v(69)
    VERIFIC_DFFRS i948 (.d(n354), .clk(clk), .s(1'b0), .r(rst), .q(m1_select[1]));   // memory_op.v(69)
    VERIFIC_DFFRS i949 (.d(n355), .clk(clk), .s(1'b0), .r(rst), .q(m1_select[0]));   // memory_op.v(69)
    VERIFIC_DFFRS i950 (.d(n552), .clk(clk), .s(1'b0), .r(rst), .q(m2_select[2]));   // memory_op.v(69)
    VERIFIC_DFFRS i951 (.d(n553), .clk(clk), .s(1'b0), .r(rst), .q(m2_select[1]));   // memory_op.v(69)
    VERIFIC_DFFRS i952 (.d(n554), .clk(clk), .s(1'b0), .r(rst), .q(m2_select[0]));   // memory_op.v(69)
    VERIFIC_DFFRS i953 (.d(r1[31]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[31]));   // memory_op.v(69)
    VERIFIC_DFFRS i954 (.d(r1[30]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[30]));   // memory_op.v(69)
    VERIFIC_DFFRS i955 (.d(r1[29]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[29]));   // memory_op.v(69)
    VERIFIC_DFFRS i956 (.d(r1[28]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[28]));   // memory_op.v(69)
    VERIFIC_DFFRS i957 (.d(r1[27]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[27]));   // memory_op.v(69)
    VERIFIC_DFFRS i958 (.d(r1[26]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[26]));   // memory_op.v(69)
    VERIFIC_DFFRS i959 (.d(r1[25]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[25]));   // memory_op.v(69)
    VERIFIC_DFFRS i960 (.d(r1[24]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[24]));   // memory_op.v(69)
    VERIFIC_DFFRS i961 (.d(r1[23]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[23]));   // memory_op.v(69)
    VERIFIC_DFFRS i962 (.d(r1[22]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[22]));   // memory_op.v(69)
    VERIFIC_DFFRS i963 (.d(r1[21]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[21]));   // memory_op.v(69)
    VERIFIC_DFFRS i964 (.d(r1[20]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[20]));   // memory_op.v(69)
    VERIFIC_DFFRS i965 (.d(r1[19]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[19]));   // memory_op.v(69)
    VERIFIC_DFFRS i966 (.d(r1[18]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[18]));   // memory_op.v(69)
    VERIFIC_DFFRS i967 (.d(r1[17]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[17]));   // memory_op.v(69)
    VERIFIC_DFFRS i968 (.d(r1[16]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[16]));   // memory_op.v(69)
    VERIFIC_DFFRS i969 (.d(r1[15]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[15]));   // memory_op.v(69)
    VERIFIC_DFFRS i970 (.d(r1[14]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[14]));   // memory_op.v(69)
    VERIFIC_DFFRS i971 (.d(r1[13]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[13]));   // memory_op.v(69)
    VERIFIC_DFFRS i972 (.d(r1[12]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[12]));   // memory_op.v(69)
    VERIFIC_DFFRS i973 (.d(r1[11]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[11]));   // memory_op.v(69)
    VERIFIC_DFFRS i974 (.d(r1[10]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[10]));   // memory_op.v(69)
    VERIFIC_DFFRS i975 (.d(r1[9]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[9]));   // memory_op.v(69)
    VERIFIC_DFFRS i976 (.d(r1[8]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[8]));   // memory_op.v(69)
    VERIFIC_DFFRS i977 (.d(r1[7]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[7]));   // memory_op.v(69)
    VERIFIC_DFFRS i978 (.d(r1[6]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[6]));   // memory_op.v(69)
    VERIFIC_DFFRS i979 (.d(r1[5]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[5]));   // memory_op.v(69)
    VERIFIC_DFFRS i980 (.d(r1[4]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[4]));   // memory_op.v(69)
    VERIFIC_DFFRS i981 (.d(r1[3]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[3]));   // memory_op.v(69)
    VERIFIC_DFFRS i982 (.d(r1[2]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[2]));   // memory_op.v(69)
    VERIFIC_DFFRS i983 (.d(r1[1]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[1]));   // memory_op.v(69)
    VERIFIC_DFFRS i984 (.d(r1[0]), .clk(clk), .s(1'b0), .r(rst), .q(r1_inner[0]));   // memory_op.v(69)
    VERIFIC_DFFRS i985 (.d(r2[31]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[31]));   // memory_op.v(69)
    VERIFIC_DFFRS i986 (.d(r2[30]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[30]));   // memory_op.v(69)
    VERIFIC_DFFRS i987 (.d(r2[29]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[29]));   // memory_op.v(69)
    VERIFIC_DFFRS i988 (.d(r2[28]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[28]));   // memory_op.v(69)
    VERIFIC_DFFRS i989 (.d(r2[27]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[27]));   // memory_op.v(69)
    VERIFIC_DFFRS i990 (.d(r2[26]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[26]));   // memory_op.v(69)
    VERIFIC_DFFRS i991 (.d(r2[25]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[25]));   // memory_op.v(69)
    VERIFIC_DFFRS i992 (.d(r2[24]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[24]));   // memory_op.v(69)
    VERIFIC_DFFRS i993 (.d(r2[23]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[23]));   // memory_op.v(69)
    VERIFIC_DFFRS i994 (.d(r2[22]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[22]));   // memory_op.v(69)
    VERIFIC_DFFRS i995 (.d(r2[21]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[21]));   // memory_op.v(69)
    VERIFIC_DFFRS i996 (.d(r2[20]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[20]));   // memory_op.v(69)
    VERIFIC_DFFRS i997 (.d(r2[19]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[19]));   // memory_op.v(69)
    VERIFIC_DFFRS i998 (.d(r2[18]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[18]));   // memory_op.v(69)
    VERIFIC_DFFRS i999 (.d(r2[17]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[17]));   // memory_op.v(69)
    VERIFIC_DFFRS i1000 (.d(r2[16]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[16]));   // memory_op.v(69)
    VERIFIC_DFFRS i1001 (.d(r2[15]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[15]));   // memory_op.v(69)
    VERIFIC_DFFRS i1002 (.d(r2[14]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[14]));   // memory_op.v(69)
    VERIFIC_DFFRS i1003 (.d(r2[13]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[13]));   // memory_op.v(69)
    VERIFIC_DFFRS i1004 (.d(r2[12]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[12]));   // memory_op.v(69)
    VERIFIC_DFFRS i1005 (.d(r2[11]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[11]));   // memory_op.v(69)
    VERIFIC_DFFRS i1006 (.d(r2[10]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[10]));   // memory_op.v(69)
    VERIFIC_DFFRS i1007 (.d(r2[9]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[9]));   // memory_op.v(69)
    VERIFIC_DFFRS i1008 (.d(r2[8]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[8]));   // memory_op.v(69)
    VERIFIC_DFFRS i1009 (.d(r2[7]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[7]));   // memory_op.v(69)
    VERIFIC_DFFRS i1010 (.d(r2[6]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[6]));   // memory_op.v(69)
    VERIFIC_DFFRS i1011 (.d(r2[5]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[5]));   // memory_op.v(69)
    VERIFIC_DFFRS i1012 (.d(r2[4]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[4]));   // memory_op.v(69)
    VERIFIC_DFFRS i1013 (.d(r2[3]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[3]));   // memory_op.v(69)
    VERIFIC_DFFRS i1014 (.d(r2[2]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[2]));   // memory_op.v(69)
    VERIFIC_DFFRS i1015 (.d(r2[1]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[1]));   // memory_op.v(69)
    VERIFIC_DFFRS i1016 (.d(r2[0]), .clk(clk), .s(1'b0), .r(rst), .q(r2_inner[0]));   // memory_op.v(69)
    VERIFIC_DFFRS i751 (.d(n685), .clk(clk), .s(1'b0), .r(rst), .q(ram_w_addr[31]));   // memory_op.v(69)
    
endmodule

//
// Verific Verilog Description of module memory_op_stage_passthrough
//

module memory_op_stage_passthrough (q_a1, q_a2, q_op, q_proceed, a1, 
            a2, op, proceed, clk, rst);   // memory_op.v(3)
    output [4:0]q_a1;   // memory_op.v(10)
    output [4:0]q_a2;   // memory_op.v(10)
    output [3:0]q_op;   // memory_op.v(11)
    output q_proceed;   // memory_op.v(12)
    input [4:0]a1;   // memory_op.v(4)
    input [4:0]a2;   // memory_op.v(4)
    input [3:0]op;   // memory_op.v(5)
    input proceed;   // memory_op.v(6)
    input clk;   // memory_op.v(8)
    input rst;   // memory_op.v(8)
    
    
    VERIFIC_DFFRS i6 (.d(a1[3]), .clk(clk), .s(1'b0), .r(rst), .q(q_a1[3]));   // memory_op.v(20)
    VERIFIC_DFFRS i7 (.d(a1[2]), .clk(clk), .s(1'b0), .r(rst), .q(q_a1[2]));   // memory_op.v(20)
    VERIFIC_DFFRS i8 (.d(a1[1]), .clk(clk), .s(1'b0), .r(rst), .q(q_a1[1]));   // memory_op.v(20)
    VERIFIC_DFFRS i9 (.d(a1[0]), .clk(clk), .s(1'b0), .r(rst), .q(q_a1[0]));   // memory_op.v(20)
    VERIFIC_DFFRS i10 (.d(a2[4]), .clk(clk), .s(1'b0), .r(rst), .q(q_a2[4]));   // memory_op.v(20)
    VERIFIC_DFFRS i11 (.d(a2[3]), .clk(clk), .s(1'b0), .r(rst), .q(q_a2[3]));   // memory_op.v(20)
    VERIFIC_DFFRS i12 (.d(a2[2]), .clk(clk), .s(1'b0), .r(rst), .q(q_a2[2]));   // memory_op.v(20)
    VERIFIC_DFFRS i13 (.d(a2[1]), .clk(clk), .s(1'b0), .r(rst), .q(q_a2[1]));   // memory_op.v(20)
    VERIFIC_DFFRS i14 (.d(a2[0]), .clk(clk), .s(1'b0), .r(rst), .q(q_a2[0]));   // memory_op.v(20)
    VERIFIC_DFFRS i15 (.d(op[3]), .clk(clk), .s(1'b0), .r(rst), .q(q_op[3]));   // memory_op.v(20)
    VERIFIC_DFFRS i16 (.d(op[2]), .clk(clk), .s(1'b0), .r(rst), .q(q_op[2]));   // memory_op.v(20)
    VERIFIC_DFFRS i17 (.d(op[1]), .clk(clk), .s(1'b0), .r(rst), .q(q_op[1]));   // memory_op.v(20)
    VERIFIC_DFFRS i18 (.d(op[0]), .clk(clk), .s(1'b0), .r(rst), .q(q_op[0]));   // memory_op.v(20)
    VERIFIC_DFFRS i19 (.d(proceed), .clk(clk), .s(1'b0), .r(rst), .q(q_proceed));   // memory_op.v(20)
    VERIFIC_DFFRS i5 (.d(a1[4]), .clk(clk), .s(1'b0), .r(rst), .q(q_a1[4]));   // memory_op.v(20)
    
endmodule

//
// Verific Verilog Description of module register_wb
//

module register_wb (write, wr1, wr2, wa1, wa2, r1, r2, a1, a2, 
            op, proceed, clk, rst);   // register_wb.v(3)
    output [1:0]write;   // register_wb.v(15)
    output [31:0]wr1;   // register_wb.v(13)
    output [31:0]wr2;   // register_wb.v(13)
    output [4:0]wa1;   // register_wb.v(14)
    output [4:0]wa2;   // register_wb.v(14)
    input [31:0]r1;   // register_wb.v(4)
    input [31:0]r2;   // register_wb.v(4)
    input [4:0]a1;   // register_wb.v(5)
    input [4:0]a2;   // register_wb.v(5)
    input [3:0]op;   // register_wb.v(7)
    input proceed;   // register_wb.v(9)
    input clk;   // register_wb.v(11)
    input rst;   // register_wb.v(11)
    
    wire [3:0]inner_op;   // register_wb.v(17)
    
    wire n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
        n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, 
        n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
        n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, 
        n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
        n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
        n79, n80, n81, n82, n83, n84;
    
    assign inner_op[3] = proceed ? op[3] : 1'b0;   // register_wb.v(19)
    assign inner_op[2] = proceed ? op[2] : 1'b0;   // register_wb.v(19)
    assign inner_op[1] = proceed ? op[1] : 1'b0;   // register_wb.v(19)
    assign inner_op[0] = proceed ? op[0] : 1'b0;   // register_wb.v(19)
    Mux_4u_16u Mux_8 (.sel({inner_op}), .data({wr1[31], wr1[31], wr1[31], 
            wr1[31], wr1[31], wr1[31], wr1[31], r1[31], r1[31], 
            r2[31], r2[31], r2[31], r1[31], r1[31], r1[31], wr1[31]}), 
            .o(n9));   // register_wb.v(29)
    Mux_4u_16u Mux_9 (.sel({inner_op}), .data({wr1[30], wr1[30], wr1[30], 
            wr1[30], wr1[30], wr1[30], wr1[30], r1[30], r1[30], 
            r2[30], r2[30], r2[30], r1[30], r1[30], r1[30], wr1[30]}), 
            .o(n10));   // register_wb.v(29)
    Mux_4u_16u Mux_10 (.sel({inner_op}), .data({wr1[29], wr1[29], wr1[29], 
            wr1[29], wr1[29], wr1[29], wr1[29], r1[29], r1[29], 
            r2[29], r2[29], r2[29], r1[29], r1[29], r1[29], wr1[29]}), 
            .o(n11));   // register_wb.v(29)
    Mux_4u_16u Mux_11 (.sel({inner_op}), .data({wr1[28], wr1[28], wr1[28], 
            wr1[28], wr1[28], wr1[28], wr1[28], r1[28], r1[28], 
            r2[28], r2[28], r2[28], r1[28], r1[28], r1[28], wr1[28]}), 
            .o(n12));   // register_wb.v(29)
    Mux_4u_16u Mux_12 (.sel({inner_op}), .data({wr1[27], wr1[27], wr1[27], 
            wr1[27], wr1[27], wr1[27], wr1[27], r1[27], r1[27], 
            r2[27], r2[27], r2[27], r1[27], r1[27], r1[27], wr1[27]}), 
            .o(n13));   // register_wb.v(29)
    Mux_4u_16u Mux_13 (.sel({inner_op}), .data({wr1[26], wr1[26], wr1[26], 
            wr1[26], wr1[26], wr1[26], wr1[26], r1[26], r1[26], 
            r2[26], r2[26], r2[26], r1[26], r1[26], r1[26], wr1[26]}), 
            .o(n14));   // register_wb.v(29)
    Mux_4u_16u Mux_14 (.sel({inner_op}), .data({wr1[25], wr1[25], wr1[25], 
            wr1[25], wr1[25], wr1[25], wr1[25], r1[25], r1[25], 
            r2[25], r2[25], r2[25], r1[25], r1[25], r1[25], wr1[25]}), 
            .o(n15));   // register_wb.v(29)
    Mux_4u_16u Mux_15 (.sel({inner_op}), .data({wr1[24], wr1[24], wr1[24], 
            wr1[24], wr1[24], wr1[24], wr1[24], r1[24], r1[24], 
            r2[24], r2[24], r2[24], r1[24], r1[24], r1[24], wr1[24]}), 
            .o(n16));   // register_wb.v(29)
    Mux_4u_16u Mux_16 (.sel({inner_op}), .data({wr1[23], wr1[23], wr1[23], 
            wr1[23], wr1[23], wr1[23], wr1[23], r1[23], r1[23], 
            r2[23], r2[23], r2[23], r1[23], r1[23], r1[23], wr1[23]}), 
            .o(n17));   // register_wb.v(29)
    Mux_4u_16u Mux_17 (.sel({inner_op}), .data({wr1[22], wr1[22], wr1[22], 
            wr1[22], wr1[22], wr1[22], wr1[22], r1[22], r1[22], 
            r2[22], r2[22], r2[22], r1[22], r1[22], r1[22], wr1[22]}), 
            .o(n18));   // register_wb.v(29)
    Mux_4u_16u Mux_18 (.sel({inner_op}), .data({wr1[21], wr1[21], wr1[21], 
            wr1[21], wr1[21], wr1[21], wr1[21], r1[21], r1[21], 
            r2[21], r2[21], r2[21], r1[21], r1[21], r1[21], wr1[21]}), 
            .o(n19));   // register_wb.v(29)
    Mux_4u_16u Mux_19 (.sel({inner_op}), .data({wr1[20], wr1[20], wr1[20], 
            wr1[20], wr1[20], wr1[20], wr1[20], r1[20], r1[20], 
            r2[20], r2[20], r2[20], r1[20], r1[20], r1[20], wr1[20]}), 
            .o(n20));   // register_wb.v(29)
    Mux_4u_16u Mux_20 (.sel({inner_op}), .data({wr1[19], wr1[19], wr1[19], 
            wr1[19], wr1[19], wr1[19], wr1[19], r1[19], r1[19], 
            r2[19], r2[19], r2[19], r1[19], r1[19], r1[19], wr1[19]}), 
            .o(n21));   // register_wb.v(29)
    Mux_4u_16u Mux_21 (.sel({inner_op}), .data({wr1[18], wr1[18], wr1[18], 
            wr1[18], wr1[18], wr1[18], wr1[18], r1[18], r1[18], 
            r2[18], r2[18], r2[18], r1[18], r1[18], r1[18], wr1[18]}), 
            .o(n22));   // register_wb.v(29)
    Mux_4u_16u Mux_22 (.sel({inner_op}), .data({wr1[17], wr1[17], wr1[17], 
            wr1[17], wr1[17], wr1[17], wr1[17], r1[17], r1[17], 
            r2[17], r2[17], r2[17], r1[17], r1[17], r1[17], wr1[17]}), 
            .o(n23));   // register_wb.v(29)
    Mux_4u_16u Mux_23 (.sel({inner_op}), .data({wr1[16], wr1[16], wr1[16], 
            wr1[16], wr1[16], wr1[16], wr1[16], r1[16], r1[16], 
            r2[16], r2[16], r2[16], r1[16], r1[16], r1[16], wr1[16]}), 
            .o(n24));   // register_wb.v(29)
    Mux_4u_16u Mux_24 (.sel({inner_op}), .data({wr1[15], wr1[15], wr1[15], 
            wr1[15], wr1[15], wr1[15], wr1[15], r1[15], r1[15], 
            r2[15], r2[15], r2[15], r1[15], r1[15], r1[15], wr1[15]}), 
            .o(n25));   // register_wb.v(29)
    Mux_4u_16u Mux_25 (.sel({inner_op}), .data({wr1[14], wr1[14], wr1[14], 
            wr1[14], wr1[14], wr1[14], wr1[14], r1[14], r1[14], 
            r2[14], r2[14], r2[14], r1[14], r1[14], r1[14], wr1[14]}), 
            .o(n26));   // register_wb.v(29)
    Mux_4u_16u Mux_26 (.sel({inner_op}), .data({wr1[13], wr1[13], wr1[13], 
            wr1[13], wr1[13], wr1[13], wr1[13], r1[13], r1[13], 
            r2[13], r2[13], r2[13], r1[13], r1[13], r1[13], wr1[13]}), 
            .o(n27));   // register_wb.v(29)
    Mux_4u_16u Mux_27 (.sel({inner_op}), .data({wr1[12], wr1[12], wr1[12], 
            wr1[12], wr1[12], wr1[12], wr1[12], r1[12], r1[12], 
            r2[12], r2[12], r2[12], r1[12], r1[12], r1[12], wr1[12]}), 
            .o(n28));   // register_wb.v(29)
    Mux_4u_16u Mux_28 (.sel({inner_op}), .data({wr1[11], wr1[11], wr1[11], 
            wr1[11], wr1[11], wr1[11], wr1[11], r1[11], r1[11], 
            r2[11], r2[11], r2[11], r1[11], r1[11], r1[11], wr1[11]}), 
            .o(n29));   // register_wb.v(29)
    Mux_4u_16u Mux_29 (.sel({inner_op}), .data({wr1[10], wr1[10], wr1[10], 
            wr1[10], wr1[10], wr1[10], wr1[10], r1[10], r1[10], 
            r2[10], r2[10], r2[10], r1[10], r1[10], r1[10], wr1[10]}), 
            .o(n30));   // register_wb.v(29)
    Mux_4u_16u Mux_30 (.sel({inner_op}), .data({wr1[9], wr1[9], wr1[9], 
            wr1[9], wr1[9], wr1[9], wr1[9], r1[9], r1[9], r2[9], 
            r2[9], r2[9], r1[9], r1[9], r1[9], wr1[9]}), .o(n31));   // register_wb.v(29)
    Mux_4u_16u Mux_31 (.sel({inner_op}), .data({wr1[8], wr1[8], wr1[8], 
            wr1[8], wr1[8], wr1[8], wr1[8], r1[8], r1[8], r2[8], 
            r2[8], r2[8], r1[8], r1[8], r1[8], wr1[8]}), .o(n32));   // register_wb.v(29)
    Mux_4u_16u Mux_32 (.sel({inner_op}), .data({wr1[7], wr1[7], wr1[7], 
            wr1[7], wr1[7], wr1[7], wr1[7], r1[7], r1[7], r2[7], 
            r2[7], r2[7], r1[7], r1[7], r1[7], wr1[7]}), .o(n33));   // register_wb.v(29)
    Mux_4u_16u Mux_33 (.sel({inner_op}), .data({wr1[6], wr1[6], wr1[6], 
            wr1[6], wr1[6], wr1[6], wr1[6], r1[6], r1[6], r2[6], 
            r2[6], r2[6], r1[6], r1[6], r1[6], wr1[6]}), .o(n34));   // register_wb.v(29)
    Mux_4u_16u Mux_34 (.sel({inner_op}), .data({wr1[5], wr1[5], wr1[5], 
            wr1[5], wr1[5], wr1[5], wr1[5], r1[5], r1[5], r2[5], 
            r2[5], r2[5], r1[5], r1[5], r1[5], wr1[5]}), .o(n35));   // register_wb.v(29)
    Mux_4u_16u Mux_35 (.sel({inner_op}), .data({wr1[4], wr1[4], wr1[4], 
            wr1[4], wr1[4], wr1[4], wr1[4], r1[4], r1[4], r2[4], 
            r2[4], r2[4], r1[4], r1[4], r1[4], wr1[4]}), .o(n36));   // register_wb.v(29)
    Mux_4u_16u Mux_36 (.sel({inner_op}), .data({wr1[3], wr1[3], wr1[3], 
            wr1[3], wr1[3], wr1[3], wr1[3], r1[3], r1[3], r2[3], 
            r2[3], r2[3], r1[3], r1[3], r1[3], wr1[3]}), .o(n37));   // register_wb.v(29)
    Mux_4u_16u Mux_37 (.sel({inner_op}), .data({wr1[2], wr1[2], wr1[2], 
            wr1[2], wr1[2], wr1[2], wr1[2], r1[2], r1[2], r2[2], 
            r2[2], r2[2], r1[2], r1[2], r1[2], wr1[2]}), .o(n38));   // register_wb.v(29)
    Mux_4u_16u Mux_38 (.sel({inner_op}), .data({wr1[1], wr1[1], wr1[1], 
            wr1[1], wr1[1], wr1[1], wr1[1], r1[1], r1[1], r2[1], 
            r2[1], r2[1], r1[1], r1[1], r1[1], wr1[1]}), .o(n39));   // register_wb.v(29)
    Mux_4u_16u Mux_39 (.sel({inner_op}), .data({wr1[0], wr1[0], wr1[0], 
            wr1[0], wr1[0], wr1[0], wr1[0], r1[0], r1[0], r2[0], 
            r2[0], r2[0], r1[0], r1[0], r1[0], wr1[0]}), .o(n40));   // register_wb.v(29)
    Mux_4u_16u Mux_40 (.sel({inner_op}), .data({wr2[31], wr2[31], wr2[31], 
            wr2[31], wr2[31], wr2[31], wr2[31], r2[31], r2[31], 
            wr2[31], wr2[31], wr2[31], wr2[31], wr2[31], wr2[31], 
            wr2[31]}), .o(n41));   // register_wb.v(29)
    Mux_4u_16u Mux_41 (.sel({inner_op}), .data({wr2[30], wr2[30], wr2[30], 
            wr2[30], wr2[30], wr2[30], wr2[30], r2[30], r2[30], 
            wr2[30], wr2[30], wr2[30], wr2[30], wr2[30], wr2[30], 
            wr2[30]}), .o(n42));   // register_wb.v(29)
    Mux_4u_16u Mux_42 (.sel({inner_op}), .data({wr2[29], wr2[29], wr2[29], 
            wr2[29], wr2[29], wr2[29], wr2[29], r2[29], r2[29], 
            wr2[29], wr2[29], wr2[29], wr2[29], wr2[29], wr2[29], 
            wr2[29]}), .o(n43));   // register_wb.v(29)
    Mux_4u_16u Mux_43 (.sel({inner_op}), .data({wr2[28], wr2[28], wr2[28], 
            wr2[28], wr2[28], wr2[28], wr2[28], r2[28], r2[28], 
            wr2[28], wr2[28], wr2[28], wr2[28], wr2[28], wr2[28], 
            wr2[28]}), .o(n44));   // register_wb.v(29)
    Mux_4u_16u Mux_44 (.sel({inner_op}), .data({wr2[27], wr2[27], wr2[27], 
            wr2[27], wr2[27], wr2[27], wr2[27], r2[27], r2[27], 
            wr2[27], wr2[27], wr2[27], wr2[27], wr2[27], wr2[27], 
            wr2[27]}), .o(n45));   // register_wb.v(29)
    Mux_4u_16u Mux_45 (.sel({inner_op}), .data({wr2[26], wr2[26], wr2[26], 
            wr2[26], wr2[26], wr2[26], wr2[26], r2[26], r2[26], 
            wr2[26], wr2[26], wr2[26], wr2[26], wr2[26], wr2[26], 
            wr2[26]}), .o(n46));   // register_wb.v(29)
    Mux_4u_16u Mux_46 (.sel({inner_op}), .data({wr2[25], wr2[25], wr2[25], 
            wr2[25], wr2[25], wr2[25], wr2[25], r2[25], r2[25], 
            wr2[25], wr2[25], wr2[25], wr2[25], wr2[25], wr2[25], 
            wr2[25]}), .o(n47));   // register_wb.v(29)
    Mux_4u_16u Mux_47 (.sel({inner_op}), .data({wr2[24], wr2[24], wr2[24], 
            wr2[24], wr2[24], wr2[24], wr2[24], r2[24], r2[24], 
            wr2[24], wr2[24], wr2[24], wr2[24], wr2[24], wr2[24], 
            wr2[24]}), .o(n48));   // register_wb.v(29)
    Mux_4u_16u Mux_48 (.sel({inner_op}), .data({wr2[23], wr2[23], wr2[23], 
            wr2[23], wr2[23], wr2[23], wr2[23], r2[23], r2[23], 
            wr2[23], wr2[23], wr2[23], wr2[23], wr2[23], wr2[23], 
            wr2[23]}), .o(n49));   // register_wb.v(29)
    Mux_4u_16u Mux_49 (.sel({inner_op}), .data({wr2[22], wr2[22], wr2[22], 
            wr2[22], wr2[22], wr2[22], wr2[22], r2[22], r2[22], 
            wr2[22], wr2[22], wr2[22], wr2[22], wr2[22], wr2[22], 
            wr2[22]}), .o(n50));   // register_wb.v(29)
    Mux_4u_16u Mux_50 (.sel({inner_op}), .data({wr2[21], wr2[21], wr2[21], 
            wr2[21], wr2[21], wr2[21], wr2[21], r2[21], r2[21], 
            wr2[21], wr2[21], wr2[21], wr2[21], wr2[21], wr2[21], 
            wr2[21]}), .o(n51));   // register_wb.v(29)
    Mux_4u_16u Mux_51 (.sel({inner_op}), .data({wr2[20], wr2[20], wr2[20], 
            wr2[20], wr2[20], wr2[20], wr2[20], r2[20], r2[20], 
            wr2[20], wr2[20], wr2[20], wr2[20], wr2[20], wr2[20], 
            wr2[20]}), .o(n52));   // register_wb.v(29)
    Mux_4u_16u Mux_52 (.sel({inner_op}), .data({wr2[19], wr2[19], wr2[19], 
            wr2[19], wr2[19], wr2[19], wr2[19], r2[19], r2[19], 
            wr2[19], wr2[19], wr2[19], wr2[19], wr2[19], wr2[19], 
            wr2[19]}), .o(n53));   // register_wb.v(29)
    Mux_4u_16u Mux_53 (.sel({inner_op}), .data({wr2[18], wr2[18], wr2[18], 
            wr2[18], wr2[18], wr2[18], wr2[18], r2[18], r2[18], 
            wr2[18], wr2[18], wr2[18], wr2[18], wr2[18], wr2[18], 
            wr2[18]}), .o(n54));   // register_wb.v(29)
    Mux_4u_16u Mux_54 (.sel({inner_op}), .data({wr2[17], wr2[17], wr2[17], 
            wr2[17], wr2[17], wr2[17], wr2[17], r2[17], r2[17], 
            wr2[17], wr2[17], wr2[17], wr2[17], wr2[17], wr2[17], 
            wr2[17]}), .o(n55));   // register_wb.v(29)
    Mux_4u_16u Mux_55 (.sel({inner_op}), .data({wr2[16], wr2[16], wr2[16], 
            wr2[16], wr2[16], wr2[16], wr2[16], r2[16], r2[16], 
            wr2[16], wr2[16], wr2[16], wr2[16], wr2[16], wr2[16], 
            wr2[16]}), .o(n56));   // register_wb.v(29)
    Mux_4u_16u Mux_56 (.sel({inner_op}), .data({wr2[15], wr2[15], wr2[15], 
            wr2[15], wr2[15], wr2[15], wr2[15], r2[15], r2[15], 
            wr2[15], wr2[15], wr2[15], wr2[15], wr2[15], wr2[15], 
            wr2[15]}), .o(n57));   // register_wb.v(29)
    Mux_4u_16u Mux_57 (.sel({inner_op}), .data({wr2[14], wr2[14], wr2[14], 
            wr2[14], wr2[14], wr2[14], wr2[14], r2[14], r2[14], 
            wr2[14], wr2[14], wr2[14], wr2[14], wr2[14], wr2[14], 
            wr2[14]}), .o(n58));   // register_wb.v(29)
    Mux_4u_16u Mux_58 (.sel({inner_op}), .data({wr2[13], wr2[13], wr2[13], 
            wr2[13], wr2[13], wr2[13], wr2[13], r2[13], r2[13], 
            wr2[13], wr2[13], wr2[13], wr2[13], wr2[13], wr2[13], 
            wr2[13]}), .o(n59));   // register_wb.v(29)
    Mux_4u_16u Mux_59 (.sel({inner_op}), .data({wr2[12], wr2[12], wr2[12], 
            wr2[12], wr2[12], wr2[12], wr2[12], r2[12], r2[12], 
            wr2[12], wr2[12], wr2[12], wr2[12], wr2[12], wr2[12], 
            wr2[12]}), .o(n60));   // register_wb.v(29)
    Mux_4u_16u Mux_60 (.sel({inner_op}), .data({wr2[11], wr2[11], wr2[11], 
            wr2[11], wr2[11], wr2[11], wr2[11], r2[11], r2[11], 
            wr2[11], wr2[11], wr2[11], wr2[11], wr2[11], wr2[11], 
            wr2[11]}), .o(n61));   // register_wb.v(29)
    Mux_4u_16u Mux_61 (.sel({inner_op}), .data({wr2[10], wr2[10], wr2[10], 
            wr2[10], wr2[10], wr2[10], wr2[10], r2[10], r2[10], 
            wr2[10], wr2[10], wr2[10], wr2[10], wr2[10], wr2[10], 
            wr2[10]}), .o(n62));   // register_wb.v(29)
    Mux_4u_16u Mux_62 (.sel({inner_op}), .data({wr2[9], wr2[9], wr2[9], 
            wr2[9], wr2[9], wr2[9], wr2[9], r2[9], r2[9], wr2[9], 
            wr2[9], wr2[9], wr2[9], wr2[9], wr2[9], wr2[9]}), .o(n63));   // register_wb.v(29)
    Mux_4u_16u Mux_63 (.sel({inner_op}), .data({wr2[8], wr2[8], wr2[8], 
            wr2[8], wr2[8], wr2[8], wr2[8], r2[8], r2[8], wr2[8], 
            wr2[8], wr2[8], wr2[8], wr2[8], wr2[8], wr2[8]}), .o(n64));   // register_wb.v(29)
    Mux_4u_16u Mux_64 (.sel({inner_op}), .data({wr2[7], wr2[7], wr2[7], 
            wr2[7], wr2[7], wr2[7], wr2[7], r2[7], r2[7], wr2[7], 
            wr2[7], wr2[7], wr2[7], wr2[7], wr2[7], wr2[7]}), .o(n65));   // register_wb.v(29)
    Mux_4u_16u Mux_65 (.sel({inner_op}), .data({wr2[6], wr2[6], wr2[6], 
            wr2[6], wr2[6], wr2[6], wr2[6], r2[6], r2[6], wr2[6], 
            wr2[6], wr2[6], wr2[6], wr2[6], wr2[6], wr2[6]}), .o(n66));   // register_wb.v(29)
    Mux_4u_16u Mux_66 (.sel({inner_op}), .data({wr2[5], wr2[5], wr2[5], 
            wr2[5], wr2[5], wr2[5], wr2[5], r2[5], r2[5], wr2[5], 
            wr2[5], wr2[5], wr2[5], wr2[5], wr2[5], wr2[5]}), .o(n67));   // register_wb.v(29)
    Mux_4u_16u Mux_67 (.sel({inner_op}), .data({wr2[4], wr2[4], wr2[4], 
            wr2[4], wr2[4], wr2[4], wr2[4], r2[4], r2[4], wr2[4], 
            wr2[4], wr2[4], wr2[4], wr2[4], wr2[4], wr2[4]}), .o(n68));   // register_wb.v(29)
    Mux_4u_16u Mux_68 (.sel({inner_op}), .data({wr2[3], wr2[3], wr2[3], 
            wr2[3], wr2[3], wr2[3], wr2[3], r2[3], r2[3], wr2[3], 
            wr2[3], wr2[3], wr2[3], wr2[3], wr2[3], wr2[3]}), .o(n69));   // register_wb.v(29)
    Mux_4u_16u Mux_69 (.sel({inner_op}), .data({wr2[2], wr2[2], wr2[2], 
            wr2[2], wr2[2], wr2[2], wr2[2], r2[2], r2[2], wr2[2], 
            wr2[2], wr2[2], wr2[2], wr2[2], wr2[2], wr2[2]}), .o(n70));   // register_wb.v(29)
    Mux_4u_16u Mux_70 (.sel({inner_op}), .data({wr2[1], wr2[1], wr2[1], 
            wr2[1], wr2[1], wr2[1], wr2[1], r2[1], r2[1], wr2[1], 
            wr2[1], wr2[1], wr2[1], wr2[1], wr2[1], wr2[1]}), .o(n71));   // register_wb.v(29)
    Mux_4u_16u Mux_71 (.sel({inner_op}), .data({wr2[0], wr2[0], wr2[0], 
            wr2[0], wr2[0], wr2[0], wr2[0], r2[0], r2[0], wr2[0], 
            wr2[0], wr2[0], wr2[0], wr2[0], wr2[0], wr2[0]}), .o(n72));   // register_wb.v(29)
    Mux_4u_16u Mux_72 (.sel({inner_op}), .data({wa1[4], wa1[4], wa1[4], 
            wa1[4], wa1[4], wa1[4], wa1[4], a2[4], a1[4], r1[4], 
            a2[4], a1[4], r2[4], a2[4], a1[4], wa1[4]}), .o(n73));   // register_wb.v(29)
    Mux_4u_16u Mux_73 (.sel({inner_op}), .data({wa1[3], wa1[3], wa1[3], 
            wa1[3], wa1[3], wa1[3], wa1[3], a2[3], a1[3], r1[3], 
            a2[3], a1[3], r2[3], a2[3], a1[3], wa1[3]}), .o(n74));   // register_wb.v(29)
    Mux_4u_16u Mux_74 (.sel({inner_op}), .data({wa1[2], wa1[2], wa1[2], 
            wa1[2], wa1[2], wa1[2], wa1[2], a2[2], a1[2], r1[2], 
            a2[2], a1[2], r2[2], a2[2], a1[2], wa1[2]}), .o(n75));   // register_wb.v(29)
    Mux_4u_16u Mux_75 (.sel({inner_op}), .data({wa1[1], wa1[1], wa1[1], 
            wa1[1], wa1[1], wa1[1], wa1[1], a2[1], a1[1], r1[1], 
            a2[1], a1[1], r2[1], a2[1], a1[1], wa1[1]}), .o(n76));   // register_wb.v(29)
    Mux_4u_16u Mux_76 (.sel({inner_op}), .data({wa1[0], wa1[0], wa1[0], 
            wa1[0], wa1[0], wa1[0], wa1[0], a2[0], a1[0], r1[0], 
            a2[0], a1[0], r2[0], a2[0], a1[0], wa1[0]}), .o(n77));   // register_wb.v(29)
    Mux_4u_16u Mux_77 (.sel({inner_op}), .data({wa2[4], wa2[4], wa2[4], 
            wa2[4], wa2[4], wa2[4], wa2[4], a1[4], a2[4], wa2[4], 
            wa2[4], wa2[4], wa2[4], wa2[4], wa2[4], wa2[4]}), .o(n78));   // register_wb.v(29)
    Mux_4u_16u Mux_78 (.sel({inner_op}), .data({wa2[3], wa2[3], wa2[3], 
            wa2[3], wa2[3], wa2[3], wa2[3], a1[3], a2[3], wa2[3], 
            wa2[3], wa2[3], wa2[3], wa2[3], wa2[3], wa2[3]}), .o(n79));   // register_wb.v(29)
    Mux_4u_16u Mux_79 (.sel({inner_op}), .data({wa2[2], wa2[2], wa2[2], 
            wa2[2], wa2[2], wa2[2], wa2[2], a1[2], a2[2], wa2[2], 
            wa2[2], wa2[2], wa2[2], wa2[2], wa2[2], wa2[2]}), .o(n80));   // register_wb.v(29)
    Mux_4u_16u Mux_80 (.sel({inner_op}), .data({wa2[1], wa2[1], wa2[1], 
            wa2[1], wa2[1], wa2[1], wa2[1], a1[1], a2[1], wa2[1], 
            wa2[1], wa2[1], wa2[1], wa2[1], wa2[1], wa2[1]}), .o(n81));   // register_wb.v(29)
    Mux_4u_16u Mux_81 (.sel({inner_op}), .data({wa2[0], wa2[0], wa2[0], 
            wa2[0], wa2[0], wa2[0], wa2[0], a1[0], a2[0], wa2[0], 
            wa2[0], wa2[0], wa2[0], wa2[0], wa2[0], wa2[0]}), .o(n82));   // register_wb.v(29)
    Mux_4u_16u Mux_82 (.sel({inner_op}), .data({16'b0000000110000000}), 
            .o(n83));   // register_wb.v(29)
    Mux_4u_16u Mux_83 (.sel({inner_op}), .data({16'b0000000111111110}), 
            .o(n84));   // register_wb.v(29)
    VERIFIC_DFFRS i86 (.d(n10), .clk(clk), .s(1'b0), .r(rst), .q(wr1[30]));   // register_wb.v(27)
    VERIFIC_DFFRS i87 (.d(n11), .clk(clk), .s(1'b0), .r(rst), .q(wr1[29]));   // register_wb.v(27)
    VERIFIC_DFFRS i88 (.d(n12), .clk(clk), .s(1'b0), .r(rst), .q(wr1[28]));   // register_wb.v(27)
    VERIFIC_DFFRS i89 (.d(n13), .clk(clk), .s(1'b0), .r(rst), .q(wr1[27]));   // register_wb.v(27)
    VERIFIC_DFFRS i90 (.d(n14), .clk(clk), .s(1'b0), .r(rst), .q(wr1[26]));   // register_wb.v(27)
    VERIFIC_DFFRS i91 (.d(n15), .clk(clk), .s(1'b0), .r(rst), .q(wr1[25]));   // register_wb.v(27)
    VERIFIC_DFFRS i92 (.d(n16), .clk(clk), .s(1'b0), .r(rst), .q(wr1[24]));   // register_wb.v(27)
    VERIFIC_DFFRS i93 (.d(n17), .clk(clk), .s(1'b0), .r(rst), .q(wr1[23]));   // register_wb.v(27)
    VERIFIC_DFFRS i94 (.d(n18), .clk(clk), .s(1'b0), .r(rst), .q(wr1[22]));   // register_wb.v(27)
    VERIFIC_DFFRS i95 (.d(n19), .clk(clk), .s(1'b0), .r(rst), .q(wr1[21]));   // register_wb.v(27)
    VERIFIC_DFFRS i96 (.d(n20), .clk(clk), .s(1'b0), .r(rst), .q(wr1[20]));   // register_wb.v(27)
    VERIFIC_DFFRS i97 (.d(n21), .clk(clk), .s(1'b0), .r(rst), .q(wr1[19]));   // register_wb.v(27)
    VERIFIC_DFFRS i98 (.d(n22), .clk(clk), .s(1'b0), .r(rst), .q(wr1[18]));   // register_wb.v(27)
    VERIFIC_DFFRS i99 (.d(n23), .clk(clk), .s(1'b0), .r(rst), .q(wr1[17]));   // register_wb.v(27)
    VERIFIC_DFFRS i100 (.d(n24), .clk(clk), .s(1'b0), .r(rst), .q(wr1[16]));   // register_wb.v(27)
    VERIFIC_DFFRS i101 (.d(n25), .clk(clk), .s(1'b0), .r(rst), .q(wr1[15]));   // register_wb.v(27)
    VERIFIC_DFFRS i102 (.d(n26), .clk(clk), .s(1'b0), .r(rst), .q(wr1[14]));   // register_wb.v(27)
    VERIFIC_DFFRS i103 (.d(n27), .clk(clk), .s(1'b0), .r(rst), .q(wr1[13]));   // register_wb.v(27)
    VERIFIC_DFFRS i104 (.d(n28), .clk(clk), .s(1'b0), .r(rst), .q(wr1[12]));   // register_wb.v(27)
    VERIFIC_DFFRS i105 (.d(n29), .clk(clk), .s(1'b0), .r(rst), .q(wr1[11]));   // register_wb.v(27)
    VERIFIC_DFFRS i106 (.d(n30), .clk(clk), .s(1'b0), .r(rst), .q(wr1[10]));   // register_wb.v(27)
    VERIFIC_DFFRS i107 (.d(n31), .clk(clk), .s(1'b0), .r(rst), .q(wr1[9]));   // register_wb.v(27)
    VERIFIC_DFFRS i108 (.d(n32), .clk(clk), .s(1'b0), .r(rst), .q(wr1[8]));   // register_wb.v(27)
    VERIFIC_DFFRS i109 (.d(n33), .clk(clk), .s(1'b0), .r(rst), .q(wr1[7]));   // register_wb.v(27)
    VERIFIC_DFFRS i110 (.d(n34), .clk(clk), .s(1'b0), .r(rst), .q(wr1[6]));   // register_wb.v(27)
    VERIFIC_DFFRS i111 (.d(n35), .clk(clk), .s(1'b0), .r(rst), .q(wr1[5]));   // register_wb.v(27)
    VERIFIC_DFFRS i112 (.d(n36), .clk(clk), .s(1'b0), .r(rst), .q(wr1[4]));   // register_wb.v(27)
    VERIFIC_DFFRS i113 (.d(n37), .clk(clk), .s(1'b0), .r(rst), .q(wr1[3]));   // register_wb.v(27)
    VERIFIC_DFFRS i114 (.d(n38), .clk(clk), .s(1'b0), .r(rst), .q(wr1[2]));   // register_wb.v(27)
    VERIFIC_DFFRS i115 (.d(n39), .clk(clk), .s(1'b0), .r(rst), .q(wr1[1]));   // register_wb.v(27)
    VERIFIC_DFFRS i116 (.d(n40), .clk(clk), .s(1'b0), .r(rst), .q(wr1[0]));   // register_wb.v(27)
    VERIFIC_DFFRS i117 (.d(n41), .clk(clk), .s(1'b0), .r(rst), .q(wr2[31]));   // register_wb.v(27)
    VERIFIC_DFFRS i118 (.d(n42), .clk(clk), .s(1'b0), .r(rst), .q(wr2[30]));   // register_wb.v(27)
    VERIFIC_DFFRS i119 (.d(n43), .clk(clk), .s(1'b0), .r(rst), .q(wr2[29]));   // register_wb.v(27)
    VERIFIC_DFFRS i120 (.d(n44), .clk(clk), .s(1'b0), .r(rst), .q(wr2[28]));   // register_wb.v(27)
    VERIFIC_DFFRS i121 (.d(n45), .clk(clk), .s(1'b0), .r(rst), .q(wr2[27]));   // register_wb.v(27)
    VERIFIC_DFFRS i122 (.d(n46), .clk(clk), .s(1'b0), .r(rst), .q(wr2[26]));   // register_wb.v(27)
    VERIFIC_DFFRS i123 (.d(n47), .clk(clk), .s(1'b0), .r(rst), .q(wr2[25]));   // register_wb.v(27)
    VERIFIC_DFFRS i124 (.d(n48), .clk(clk), .s(1'b0), .r(rst), .q(wr2[24]));   // register_wb.v(27)
    VERIFIC_DFFRS i125 (.d(n49), .clk(clk), .s(1'b0), .r(rst), .q(wr2[23]));   // register_wb.v(27)
    VERIFIC_DFFRS i126 (.d(n50), .clk(clk), .s(1'b0), .r(rst), .q(wr2[22]));   // register_wb.v(27)
    VERIFIC_DFFRS i127 (.d(n51), .clk(clk), .s(1'b0), .r(rst), .q(wr2[21]));   // register_wb.v(27)
    VERIFIC_DFFRS i128 (.d(n52), .clk(clk), .s(1'b0), .r(rst), .q(wr2[20]));   // register_wb.v(27)
    VERIFIC_DFFRS i129 (.d(n53), .clk(clk), .s(1'b0), .r(rst), .q(wr2[19]));   // register_wb.v(27)
    VERIFIC_DFFRS i130 (.d(n54), .clk(clk), .s(1'b0), .r(rst), .q(wr2[18]));   // register_wb.v(27)
    VERIFIC_DFFRS i131 (.d(n55), .clk(clk), .s(1'b0), .r(rst), .q(wr2[17]));   // register_wb.v(27)
    VERIFIC_DFFRS i132 (.d(n56), .clk(clk), .s(1'b0), .r(rst), .q(wr2[16]));   // register_wb.v(27)
    VERIFIC_DFFRS i133 (.d(n57), .clk(clk), .s(1'b0), .r(rst), .q(wr2[15]));   // register_wb.v(27)
    VERIFIC_DFFRS i134 (.d(n58), .clk(clk), .s(1'b0), .r(rst), .q(wr2[14]));   // register_wb.v(27)
    VERIFIC_DFFRS i135 (.d(n59), .clk(clk), .s(1'b0), .r(rst), .q(wr2[13]));   // register_wb.v(27)
    VERIFIC_DFFRS i136 (.d(n60), .clk(clk), .s(1'b0), .r(rst), .q(wr2[12]));   // register_wb.v(27)
    VERIFIC_DFFRS i137 (.d(n61), .clk(clk), .s(1'b0), .r(rst), .q(wr2[11]));   // register_wb.v(27)
    VERIFIC_DFFRS i138 (.d(n62), .clk(clk), .s(1'b0), .r(rst), .q(wr2[10]));   // register_wb.v(27)
    VERIFIC_DFFRS i139 (.d(n63), .clk(clk), .s(1'b0), .r(rst), .q(wr2[9]));   // register_wb.v(27)
    VERIFIC_DFFRS i140 (.d(n64), .clk(clk), .s(1'b0), .r(rst), .q(wr2[8]));   // register_wb.v(27)
    VERIFIC_DFFRS i141 (.d(n65), .clk(clk), .s(1'b0), .r(rst), .q(wr2[7]));   // register_wb.v(27)
    VERIFIC_DFFRS i142 (.d(n66), .clk(clk), .s(1'b0), .r(rst), .q(wr2[6]));   // register_wb.v(27)
    VERIFIC_DFFRS i143 (.d(n67), .clk(clk), .s(1'b0), .r(rst), .q(wr2[5]));   // register_wb.v(27)
    VERIFIC_DFFRS i144 (.d(n68), .clk(clk), .s(1'b0), .r(rst), .q(wr2[4]));   // register_wb.v(27)
    VERIFIC_DFFRS i145 (.d(n69), .clk(clk), .s(1'b0), .r(rst), .q(wr2[3]));   // register_wb.v(27)
    VERIFIC_DFFRS i146 (.d(n70), .clk(clk), .s(1'b0), .r(rst), .q(wr2[2]));   // register_wb.v(27)
    VERIFIC_DFFRS i147 (.d(n71), .clk(clk), .s(1'b0), .r(rst), .q(wr2[1]));   // register_wb.v(27)
    VERIFIC_DFFRS i148 (.d(n72), .clk(clk), .s(1'b0), .r(rst), .q(wr2[0]));   // register_wb.v(27)
    VERIFIC_DFFRS i149 (.d(n73), .clk(clk), .s(1'b0), .r(rst), .q(wa1[4]));   // register_wb.v(27)
    VERIFIC_DFFRS i150 (.d(n74), .clk(clk), .s(1'b0), .r(rst), .q(wa1[3]));   // register_wb.v(27)
    VERIFIC_DFFRS i151 (.d(n75), .clk(clk), .s(1'b0), .r(rst), .q(wa1[2]));   // register_wb.v(27)
    VERIFIC_DFFRS i152 (.d(n76), .clk(clk), .s(1'b0), .r(rst), .q(wa1[1]));   // register_wb.v(27)
    VERIFIC_DFFRS i153 (.d(n77), .clk(clk), .s(1'b0), .r(rst), .q(wa1[0]));   // register_wb.v(27)
    VERIFIC_DFFRS i154 (.d(n78), .clk(clk), .s(1'b0), .r(rst), .q(wa2[4]));   // register_wb.v(27)
    VERIFIC_DFFRS i155 (.d(n79), .clk(clk), .s(1'b0), .r(rst), .q(wa2[3]));   // register_wb.v(27)
    VERIFIC_DFFRS i156 (.d(n80), .clk(clk), .s(1'b0), .r(rst), .q(wa2[2]));   // register_wb.v(27)
    VERIFIC_DFFRS i157 (.d(n81), .clk(clk), .s(1'b0), .r(rst), .q(wa2[1]));   // register_wb.v(27)
    VERIFIC_DFFRS i158 (.d(n82), .clk(clk), .s(1'b0), .r(rst), .q(wa2[0]));   // register_wb.v(27)
    VERIFIC_DFFRS i159 (.d(n83), .clk(clk), .s(1'b0), .r(rst), .q(write[1]));   // register_wb.v(27)
    VERIFIC_DFFRS i160 (.d(n84), .clk(clk), .s(1'b0), .r(rst), .q(write[0]));   // register_wb.v(27)
    VERIFIC_DFFRS i85 (.d(n9), .clk(clk), .s(1'b0), .r(rst), .q(wr1[31]));   // register_wb.v(27)
    
endmodule

//
// Verific Verilog Description of module reg_hazard_checker
//

module reg_hazard_checker (ex_hazard, mem_hazard, reg_hazard, ex_r1_a, 
            ex_r2_a, ex_r_op, ex_proceed, mem_r1_a, mem_r2_a, mem_r_op, 
            mem_proceed, reg_r1_a, reg_r2_a, reg_write, dec_r1_addr, 
            dec_r2_addr, dec_r_read);   // insn_decoder.v(18)
    output ex_hazard;   // insn_decoder.v(19)
    output mem_hazard;   // insn_decoder.v(20)
    output reg_hazard;   // insn_decoder.v(21)
    input [4:0]ex_r1_a;   // insn_decoder.v(23)
    input [4:0]ex_r2_a;   // insn_decoder.v(23)
    input [3:0]ex_r_op;   // insn_decoder.v(24)
    input ex_proceed;   // insn_decoder.v(25)
    input [4:0]mem_r1_a;   // insn_decoder.v(27)
    input [4:0]mem_r2_a;   // insn_decoder.v(27)
    input [3:0]mem_r_op;   // insn_decoder.v(28)
    input mem_proceed;   // insn_decoder.v(29)
    input [4:0]reg_r1_a;   // insn_decoder.v(31)
    input [4:0]reg_r2_a;   // insn_decoder.v(31)
    input [1:0]reg_write;   // insn_decoder.v(32)
    input [4:0]dec_r1_addr;   // insn_decoder.v(34)
    input [4:0]dec_r2_addr;   // insn_decoder.v(34)
    input [1:0]dec_r_read;   // insn_decoder.v(35)
    
    wire ex_r1_op_comp;   // insn_decoder.v(40)
    wire ex_r2_op_comp;   // insn_decoder.v(41)
    wire ex_r1r2_op_comp;   // insn_decoder.v(42)
    wire ex_r1_comp;   // insn_decoder.v(44)
    wire ex_r2_comp;   // insn_decoder.v(45)
    wire ex_r1r2_comp;   // insn_decoder.v(46)
    wire ex_r2r1_comp;   // insn_decoder.v(47)
    wire ex_hazard_r1;   // insn_decoder.v(49)
    wire ex_hazard_r2;   // insn_decoder.v(50)
    wire ex_hazard_r1r2;   // insn_decoder.v(51)
    wire ex_hazard_r2r1;   // insn_decoder.v(52)
    wire mem_r1_op_comp;   // insn_decoder.v(56)
    wire mem_r2_op_comp;   // insn_decoder.v(57)
    wire mem_r1r2_op_comp;   // insn_decoder.v(58)
    wire mem_r1_comp;   // insn_decoder.v(60)
    wire mem_r2_comp;   // insn_decoder.v(61)
    wire mem_r1r2_comp;   // insn_decoder.v(62)
    wire mem_r2r1_comp;   // insn_decoder.v(63)
    wire mem_hazard_r1;   // insn_decoder.v(65)
    wire mem_hazard_r2;   // insn_decoder.v(66)
    wire mem_hazard_r1r2;   // insn_decoder.v(67)
    wire mem_hazard_r2r1;   // insn_decoder.v(68)
    wire reg_r1_comp;   // insn_decoder.v(75)
    wire reg_r2_comp;   // insn_decoder.v(76)
    wire reg_r1r2_comp;   // insn_decoder.v(77)
    wire reg_r2r1_comp;   // insn_decoder.v(78)
    wire reg_hazard_r1;   // insn_decoder.v(80)
    wire reg_hazard_r2;   // insn_decoder.v(81)
    wire reg_hazard_r1r2;   // insn_decoder.v(82)
    wire reg_hazard_r2r1;   // insn_decoder.v(83)
    
    wire n4, n5, n6, n7, n8, n11, n13, n14, n17, n18, n21, 
        n26, n27, n28, n30, n31, n32, n33, n34, n36, n37, 
        n38, n39, n40, n42, n43, n44, n45, n46, n48, n49, 
        n50, n51, n52, n54, n55, n57, n58, n61, n64, n66, 
        n67, n68, n70, n71, n72, n73, n74, n77, n79, n80, 
        n83, n84, n87, n92, n93, n94, n96, n97, n98, n99, 
        n100, n102, n103, n104, n105, n106, n108, n109, n110, 
        n111, n112, n114, n115, n116, n117, n118, n120, n121, 
        n123, n124, n127, n130, n132, n133, n134, n136, n137, 
        n138, n139, n140, n142, n143, n144, n145, n146, n148, 
        n149, n150, n151, n152, n154, n155, n156, n157, n158, 
        n160, n162, n164, n166, n168, n169;
    
    not (n4, ex_r_op[0]) ;   // insn_decoder.v(40)
    nor (n5, ex_r_op[3], ex_r_op[2], ex_r_op[1], n4) ;   // insn_decoder.v(40)
    not (n6, ex_r_op[1]) ;   // insn_decoder.v(40)
    nor (n7, ex_r_op[3], ex_r_op[2], n6, ex_r_op[0]) ;   // insn_decoder.v(40)
    or (n8, n5, n7) ;   // insn_decoder.v(40)
    nor (n11, ex_r_op[3], ex_r_op[2], n6, n4) ;   // insn_decoder.v(40)
    or (ex_r1_op_comp, n8, n11) ;   // insn_decoder.v(40)
    not (n13, ex_r_op[2]) ;   // insn_decoder.v(41)
    nor (n14, ex_r_op[3], n13, ex_r_op[1], ex_r_op[0]) ;   // insn_decoder.v(41)
    nor (n17, ex_r_op[3], n13, ex_r_op[1], n4) ;   // insn_decoder.v(41)
    or (n18, n14, n17) ;   // insn_decoder.v(41)
    nor (n21, ex_r_op[3], n13, n6, ex_r_op[0]) ;   // insn_decoder.v(41)
    or (ex_r2_op_comp, n18, n21) ;   // insn_decoder.v(41)
    nor (n26, ex_r_op[3], n13, n6, n4) ;   // insn_decoder.v(42)
    not (n27, ex_r_op[3]) ;   // insn_decoder.v(42)
    nor (n28, n27, ex_r_op[2], ex_r_op[1], ex_r_op[0]) ;   // insn_decoder.v(42)
    or (ex_r1r2_op_comp, n26, n28) ;   // insn_decoder.v(42)
    xor (n30, ex_r1_a[0], dec_r1_addr[0]) ;   // insn_decoder.v(44)
    xor (n31, ex_r1_a[1], dec_r1_addr[1]) ;   // insn_decoder.v(44)
    xor (n32, ex_r1_a[2], dec_r1_addr[2]) ;   // insn_decoder.v(44)
    xor (n33, ex_r1_a[3], dec_r1_addr[3]) ;   // insn_decoder.v(44)
    xor (n34, ex_r1_a[4], dec_r1_addr[4]) ;   // insn_decoder.v(44)
    nor (ex_r1_comp, n34, n33, n32, n31, n30) ;   // insn_decoder.v(44)
    xor (n36, ex_r2_a[0], dec_r2_addr[0]) ;   // insn_decoder.v(45)
    xor (n37, ex_r2_a[1], dec_r2_addr[1]) ;   // insn_decoder.v(45)
    xor (n38, ex_r2_a[2], dec_r2_addr[2]) ;   // insn_decoder.v(45)
    xor (n39, ex_r2_a[3], dec_r2_addr[3]) ;   // insn_decoder.v(45)
    xor (n40, ex_r2_a[4], dec_r2_addr[4]) ;   // insn_decoder.v(45)
    nor (ex_r2_comp, n40, n39, n38, n37, n36) ;   // insn_decoder.v(45)
    xor (n42, ex_r1_a[0], dec_r2_addr[0]) ;   // insn_decoder.v(46)
    xor (n43, ex_r1_a[1], dec_r2_addr[1]) ;   // insn_decoder.v(46)
    xor (n44, ex_r1_a[2], dec_r2_addr[2]) ;   // insn_decoder.v(46)
    xor (n45, ex_r1_a[3], dec_r2_addr[3]) ;   // insn_decoder.v(46)
    xor (n46, ex_r1_a[4], dec_r2_addr[4]) ;   // insn_decoder.v(46)
    nor (ex_r1r2_comp, n46, n45, n44, n43, n42) ;   // insn_decoder.v(46)
    xor (n48, ex_r2_a[0], dec_r1_addr[0]) ;   // insn_decoder.v(47)
    xor (n49, ex_r2_a[1], dec_r1_addr[1]) ;   // insn_decoder.v(47)
    xor (n50, ex_r2_a[2], dec_r1_addr[2]) ;   // insn_decoder.v(47)
    xor (n51, ex_r2_a[3], dec_r1_addr[3]) ;   // insn_decoder.v(47)
    xor (n52, ex_r2_a[4], dec_r1_addr[4]) ;   // insn_decoder.v(47)
    nor (ex_r2r1_comp, n52, n51, n50, n49, n48) ;   // insn_decoder.v(47)
    or (n54, ex_r1_op_comp, ex_r1r2_op_comp) ;   // insn_decoder.v(49)
    and (n55, n54, ex_r1_comp) ;   // insn_decoder.v(49)
    and (ex_hazard_r1, n55, dec_r_read[0]) ;   // insn_decoder.v(49)
    or (n57, ex_r2_op_comp, ex_r1r2_op_comp) ;   // insn_decoder.v(50)
    and (n58, n57, ex_r2_comp) ;   // insn_decoder.v(50)
    and (ex_hazard_r2, n58, dec_r_read[1]) ;   // insn_decoder.v(50)
    and (n61, n54, ex_r1r2_comp) ;   // insn_decoder.v(51)
    and (ex_hazard_r1r2, n61, dec_r_read[1]) ;   // insn_decoder.v(51)
    and (n64, n57, ex_r2r1_comp) ;   // insn_decoder.v(52)
    and (ex_hazard_r2r1, n64, dec_r_read[0]) ;   // insn_decoder.v(52)
    or (n66, ex_hazard_r1, ex_hazard_r2) ;   // insn_decoder.v(54)
    or (n67, n66, ex_hazard_r1r2) ;   // insn_decoder.v(54)
    or (n68, n67, ex_hazard_r2r1) ;   // insn_decoder.v(54)
    and (ex_hazard, n68, ex_proceed) ;   // insn_decoder.v(54)
    not (n70, mem_r_op[0]) ;   // insn_decoder.v(56)
    nor (n71, mem_r_op[3], mem_r_op[2], mem_r_op[1], n70) ;   // insn_decoder.v(56)
    not (n72, mem_r_op[1]) ;   // insn_decoder.v(56)
    nor (n73, mem_r_op[3], mem_r_op[2], n72, mem_r_op[0]) ;   // insn_decoder.v(56)
    or (n74, n71, n73) ;   // insn_decoder.v(56)
    nor (n77, mem_r_op[3], mem_r_op[2], n72, n70) ;   // insn_decoder.v(56)
    or (mem_r1_op_comp, n74, n77) ;   // insn_decoder.v(56)
    not (n79, mem_r_op[2]) ;   // insn_decoder.v(57)
    nor (n80, mem_r_op[3], n79, mem_r_op[1], mem_r_op[0]) ;   // insn_decoder.v(57)
    nor (n83, mem_r_op[3], n79, mem_r_op[1], n70) ;   // insn_decoder.v(57)
    or (n84, n80, n83) ;   // insn_decoder.v(57)
    nor (n87, mem_r_op[3], n79, n72, mem_r_op[0]) ;   // insn_decoder.v(57)
    or (mem_r2_op_comp, n84, n87) ;   // insn_decoder.v(57)
    nor (n92, mem_r_op[3], n79, n72, n70) ;   // insn_decoder.v(58)
    not (n93, mem_r_op[3]) ;   // insn_decoder.v(58)
    nor (n94, n93, mem_r_op[2], mem_r_op[1], mem_r_op[0]) ;   // insn_decoder.v(58)
    or (mem_r1r2_op_comp, n92, n94) ;   // insn_decoder.v(58)
    xor (n96, mem_r1_a[0], dec_r1_addr[0]) ;   // insn_decoder.v(60)
    xor (n97, mem_r1_a[1], dec_r1_addr[1]) ;   // insn_decoder.v(60)
    xor (n98, mem_r1_a[2], dec_r1_addr[2]) ;   // insn_decoder.v(60)
    xor (n99, mem_r1_a[3], dec_r1_addr[3]) ;   // insn_decoder.v(60)
    xor (n100, mem_r1_a[4], dec_r1_addr[4]) ;   // insn_decoder.v(60)
    nor (mem_r1_comp, n100, n99, n98, n97, n96) ;   // insn_decoder.v(60)
    xor (n102, mem_r2_a[0], dec_r2_addr[0]) ;   // insn_decoder.v(61)
    xor (n103, mem_r2_a[1], dec_r2_addr[1]) ;   // insn_decoder.v(61)
    xor (n104, mem_r2_a[2], dec_r2_addr[2]) ;   // insn_decoder.v(61)
    xor (n105, mem_r2_a[3], dec_r2_addr[3]) ;   // insn_decoder.v(61)
    xor (n106, mem_r2_a[4], dec_r2_addr[4]) ;   // insn_decoder.v(61)
    nor (mem_r2_comp, n106, n105, n104, n103, n102) ;   // insn_decoder.v(61)
    xor (n108, mem_r1_a[0], dec_r2_addr[0]) ;   // insn_decoder.v(62)
    xor (n109, mem_r1_a[1], dec_r2_addr[1]) ;   // insn_decoder.v(62)
    xor (n110, mem_r1_a[2], dec_r2_addr[2]) ;   // insn_decoder.v(62)
    xor (n111, mem_r1_a[3], dec_r2_addr[3]) ;   // insn_decoder.v(62)
    xor (n112, mem_r1_a[4], dec_r2_addr[4]) ;   // insn_decoder.v(62)
    nor (mem_r1r2_comp, n112, n111, n110, n109, n108) ;   // insn_decoder.v(62)
    xor (n114, mem_r2_a[0], dec_r1_addr[0]) ;   // insn_decoder.v(63)
    xor (n115, mem_r2_a[1], dec_r1_addr[1]) ;   // insn_decoder.v(63)
    xor (n116, mem_r2_a[2], dec_r1_addr[2]) ;   // insn_decoder.v(63)
    xor (n117, mem_r2_a[3], dec_r1_addr[3]) ;   // insn_decoder.v(63)
    xor (n118, mem_r2_a[4], dec_r1_addr[4]) ;   // insn_decoder.v(63)
    nor (mem_r2r1_comp, n118, n117, n116, n115, n114) ;   // insn_decoder.v(63)
    or (n120, mem_r1_op_comp, mem_r1r2_op_comp) ;   // insn_decoder.v(65)
    and (n121, n120, mem_r1_comp) ;   // insn_decoder.v(65)
    and (mem_hazard_r1, n121, dec_r_read[0]) ;   // insn_decoder.v(65)
    or (n123, mem_r2_op_comp, mem_r1r2_op_comp) ;   // insn_decoder.v(66)
    and (n124, n123, mem_r2_comp) ;   // insn_decoder.v(66)
    and (mem_hazard_r2, n124, dec_r_read[1]) ;   // insn_decoder.v(66)
    and (n127, n120, mem_r1r2_comp) ;   // insn_decoder.v(67)
    and (mem_hazard_r1r2, n127, dec_r_read[1]) ;   // insn_decoder.v(67)
    and (n130, n123, mem_r2r1_comp) ;   // insn_decoder.v(68)
    and (mem_hazard_r2r1, n130, dec_r_read[0]) ;   // insn_decoder.v(68)
    or (n132, mem_hazard_r1, mem_hazard_r2) ;   // insn_decoder.v(70)
    or (n133, n132, mem_hazard_r1r2) ;   // insn_decoder.v(70)
    or (n134, n133, mem_hazard_r2r1) ;   // insn_decoder.v(70)
    and (mem_hazard, n134, mem_proceed) ;   // insn_decoder.v(70)
    xor (n136, reg_r1_a[0], dec_r1_addr[0]) ;   // insn_decoder.v(75)
    xor (n137, reg_r1_a[1], dec_r1_addr[1]) ;   // insn_decoder.v(75)
    xor (n138, reg_r1_a[2], dec_r1_addr[2]) ;   // insn_decoder.v(75)
    xor (n139, reg_r1_a[3], dec_r1_addr[3]) ;   // insn_decoder.v(75)
    xor (n140, reg_r1_a[4], dec_r1_addr[4]) ;   // insn_decoder.v(75)
    nor (reg_r1_comp, n140, n139, n138, n137, n136) ;   // insn_decoder.v(75)
    xor (n142, reg_r2_a[0], dec_r2_addr[0]) ;   // insn_decoder.v(76)
    xor (n143, reg_r2_a[1], dec_r2_addr[1]) ;   // insn_decoder.v(76)
    xor (n144, reg_r2_a[2], dec_r2_addr[2]) ;   // insn_decoder.v(76)
    xor (n145, reg_r2_a[3], dec_r2_addr[3]) ;   // insn_decoder.v(76)
    xor (n146, reg_r2_a[4], dec_r2_addr[4]) ;   // insn_decoder.v(76)
    nor (reg_r2_comp, n146, n145, n144, n143, n142) ;   // insn_decoder.v(76)
    xor (n148, reg_r1_a[0], dec_r2_addr[0]) ;   // insn_decoder.v(77)
    xor (n149, reg_r1_a[1], dec_r2_addr[1]) ;   // insn_decoder.v(77)
    xor (n150, reg_r1_a[2], dec_r2_addr[2]) ;   // insn_decoder.v(77)
    xor (n151, reg_r1_a[3], dec_r2_addr[3]) ;   // insn_decoder.v(77)
    xor (n152, reg_r1_a[4], dec_r2_addr[4]) ;   // insn_decoder.v(77)
    nor (reg_r1r2_comp, n152, n151, n150, n149, n148) ;   // insn_decoder.v(77)
    xor (n154, reg_r2_a[0], dec_r1_addr[0]) ;   // insn_decoder.v(78)
    xor (n155, reg_r2_a[1], dec_r1_addr[1]) ;   // insn_decoder.v(78)
    xor (n156, reg_r2_a[2], dec_r1_addr[2]) ;   // insn_decoder.v(78)
    xor (n157, reg_r2_a[3], dec_r1_addr[3]) ;   // insn_decoder.v(78)
    xor (n158, reg_r2_a[4], dec_r1_addr[4]) ;   // insn_decoder.v(78)
    nor (reg_r2r1_comp, n158, n157, n156, n155, n154) ;   // insn_decoder.v(78)
    and (n160, reg_write[0], reg_r1_comp) ;   // insn_decoder.v(80)
    and (reg_hazard_r1, n160, dec_r_read[0]) ;   // insn_decoder.v(80)
    and (n162, reg_write[1], reg_r2_comp) ;   // insn_decoder.v(81)
    and (reg_hazard_r2, n162, dec_r_read[1]) ;   // insn_decoder.v(81)
    and (n164, reg_write[0], reg_r1r2_comp) ;   // insn_decoder.v(82)
    and (reg_hazard_r1r2, n164, dec_r_read[1]) ;   // insn_decoder.v(82)
    and (n166, reg_write[1], reg_r2r1_comp) ;   // insn_decoder.v(83)
    and (reg_hazard_r2r1, n166, dec_r_read[0]) ;   // insn_decoder.v(83)
    or (n168, reg_hazard_r1, reg_hazard_r2) ;   // insn_decoder.v(85)
    or (n169, n168, reg_hazard_r1r2) ;   // insn_decoder.v(85)
    or (reg_hazard, n169, reg_hazard_r2r1) ;   // insn_decoder.v(85)
    
endmodule
